`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Baig3HYrIldYL5qRvdwwMdSf0La+HeKDA6wcCFYN3GgVp5DL4jzat25zk4KWFOqT+MRI502m8fA0
Zp+CvI868A==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gAsGTvdGW2Yv3x/fbuZoBZ6DL81/fM9nG6kd5fd8TURZCo+DNNX+lRwiZtL0yiKI4mcZAbylzZ4y
a4jXbUNdghsy87GtGyL1PcVwoPBGSPQaoo7bN0CR5ENtVC7cikM5YZ6lwZ75Ckjxym3+tpTES0aJ
ovavfDx24KJv8MltNv4=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wZTGHNVSWbMoJb5A9nXjOiX6Afzz31BGrrqtPnU6jRY3JEK8eVLg1vGcTeYugU8BnjH2PCmZ/fH4
sV/2sTFS7HFFCifN8LkkaVbtMmulZC8yF56PtfHZZc61rVbCOeY4YkzYxqwuP84GrVF2RINqJ1xU
Ckzu8/Mw/iW/NBlPMAYGvntPnWlMOe29aEbb2fQSAy8SngVwlfOZQO4o9/PHhi12vEjZXC/pr4Tx
ILx2w0wwIpitm/xvh7ImdB+yOsp8LOBIW6xtXngOPT//YOzhV/mtzvuXlmel86uY4OmFnDA2colk
cOy6AqP8moAVQLd4qNda3n5PFgSh/i4IdyRVwg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tYUdeOjB2zdGhQFkEQBXD3g8osRNQGkgSNiawx6OjmC5Kk4TRW6SlIuUJNaI2IKRaTVGYELiIQPN
P49dK7Vtm3ch5MC0BIddGVCmwVk7VkrGOnw3EP6GHOqifEya1jM4ZNB1ABPFOwR6s1hYlJtLFdYJ
ZiLGBQpt7+aSoRWa0CL6nGKegUqLLMNPHSeStPvumZTzs7UU+lxs0MuwD3NGC5M/ZCDXxZXF+1dF
f4eNTFoGYq7gjml8zM88r0zXbHKbpX69jvjlEUL5jzcyWp0ae5/mSCKc04CqgxPNBv2o0hvmVO2Q
pwEfiiNAlp3gwGDoM3Hw3pdg9cx5XPN39d8MNQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mPT4AhFJbd4R7SES/GW1G2UghrfZG9KG7Jwew7gkBfFytqu+vlaBWKpAHBIQD6veLVs7PmYWoQWi
3IM7aKAkxS5m2GS1ONlgotAlcunYYXIhvU3iZyUSUJ3hNBfGiSg49OD7H6EnRMan3UvN5L5DM7Yg
Rt9224LLhImDj0UopZ0=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
scQ19a1DzcC/bww1GnRbFjlAF7M3/pkO3jtdTgiagrvmnvEq39EfKNMc88Km/beeF+e1efokRP6D
RQT6WgC4Zt25Nt8/1LzSp6MLnGVQ/wbW/od9zyg6lXk1j7CrxR7owCoGA26hqto/fBeohAkV9pJ6
S/EroO0Fy/y0pdv6hfbBE+EjRrOHiFm7FB5pQRNsB0osMmZaYJOQaGutubxIQeEIsLljSS9lR32x
4TEjPtGMMUo/cRRVtGgx73s5J+wPWalR4CMa2hheX08kZQdRJD8RwpVr4ldVdrQA7zriA5xHQOom
KH11Ut7Kxjv+LYgJ6M+rv2gZ/PPwFbvfRl3cKg==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OyEpDeJ8KK6w7Tyqv3GnJOs57gfeZ3seyKfsYCtCvlfu5FxzTKrCgUnbhdLg/ei5npcgMoyAb+Jo
8yFoPGiA43JI2oGn8NT7I72vUWa/rfdGHf+SC8fxtM41KGIPnO13xfp3Ajh/132XFXDj5YOpQALt
M47pE42FvlfrnqyWGmRBYGg7qSYEO2puEWBmxA2QNgW07twGxMu7n7ukYXjAmbodkkAML1XVd+B9
LdAAj/1QTNiIbfxyYh17N0R13rDv41yr5nE+PnmzhSekeI9mAi+DekWdYyurw5WvxtxMMQVI7Jfq
yz4tKk0faHfxpSRtwnTqSNEBbSlQy9L6VTBhhA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WlocrSfIH6PAXOhkNUeUYLueDTNKpE+nmD9Swv4croX/00MfeSXsoLW8ZAnJ8qj6tA7lMD6jFlTP
5GKRvElIf+DDiPWHfw05RmOAbtLLTfuSxVzncdSKE9cPfyfFPITG8wHqyHXUcnec7wtg4+mJmCwP
t8TUg+ZV0/fW71GeCtkK+yZG8TirR/FJJLrZvVwhkz+ui7SYbtvr2UQ872wrwPcwEycW0XlJRWKV
wAF/Ze3R9GDJgsqhSsfGeRZrzE6tZ/YyaquZMeTqJcMMrGuh6oeTzdbjR5FMyKxAfk5IUsRgKH6K
WL5lOrb1vgF/QzF/pUm1SAKSmaNxWao+DTAG1g==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PprnCfC5k/ZaA2abyUxic6Lv7c/uadKfp/cnIoehX9JA0gmQeuunNwu9D/9rCPOk1yGaw4eHdrIi
ZIVc7Y9fy8Y9F2u1sDEf7GYxr8r3qpvmgb0c9BCVlcasz8euEymGjGgG3LJTKBrU0FWXlaSC1/ek
8DxGWoQTjUknjsave1mKXVZcK08P0rLGuPD3qpiUnF+LuV3pmJ/CBA4ZV+3LWVqOwtDQ3WeRN0jF
8YjgA9INBmjXX+NHtPauCvLTWhUSNdjQ394Qu0cF4XnXV4tJ0XRe5F+BNNscr9/b9/h4U/x9WLkV
7255nZFsWz4XhTb/0zAEfi+IUWwv+vOrSCt7ZQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 98368)
`protect data_block
4gBJHPy3wv3Ip6YC0Tmqn8nSYTHoDiE/R7mj5TauEBTh+jEElE1NY3oEts/YCJJP+52VYqYm2+Bd
jNcO3qaZmacbf+XeYTKaMxPB4MHEy0inRq9/HnG90s+8k9IAXvToi/M3XSdh6e83x3LyZcO6vJIA
iYXiBvnYz2UuQxv6Zy2qqAlvlYzA42gN+Pcq38V4CTA1nk/6+JP2IvL76RgAeJSSQeiAu8VRgz6W
8A42j+m8UeDSgjWadMwW8eLhPB8yPJrfYXUG0xOR0VeQ5GWNieXcT50qgmEFENOK/b0QyJMlf44U
g2K9gEKpG04QW14idwyZELbPsOu6o7oxHRO7pZhdFxySwIILDwinhRF4QBKIJmUYPpVXPeq2DAnx
8N6yalrAWjCOjltAq80stbGWTazHhVRqvg/V6SxLbSzFUynLCj2bRdsgVvYpfu+2HaVvj3nzGamx
JR1GuVYijrsSywTYfLkMj5czC5elUhicGmiQcq6Q0U/bmcN96BycaAm5lnetVsyW0n8AqrDHlE/x
ZuFwyCkmg0prZ6lHnNX9tQz+94QNzetBdCN7lVKl8DWh3Ej0KwQzm6DpLSxCh4Tb92gKscKeJ4IP
rTHMlUH6CFNtQWksxmFK9hPoSFoBUkctMtJpARTasR/nZw6hk+XPcs2EzyKyAek54flCZ6oIHwhA
RXnF03gP4aQ22pjDXAxQCA/MSk+Zzti8AjWZWTrl83bFBwV8CU+Gr0cXv9vbWo84ByaQu1JqViPu
wTkMaHTBwdC6B/p67YemiphPRSerAkaqcQt/c+D3f/4VHiIYRojBdyPGuXVEgqGugdCJkQuoSc5v
VyC2wcW753dh8apb7BH5OeirxupGzUe9AnXrEOfu2dZM4roS5ReapYkx4BxLR99hPztWAnNWzlYV
l4iquRf1JjmjfjXuCA8oXTovt8sj31yVpgXntRd/iX9qCBP8LPfN+bCFG8FWOzV/504m03FNCVAE
BHgviXbf7XmTZzV0I3ayeDnmCCT0a0xY0HXPaOGj7DmAajjywvvyCueRMpgOXzwwldL+r1ECmCnq
tpGSTugrpqD7rY7dCMiWPXdGhiW5DR/piMn9RfKaJQx/bzBYoCAHxrxLo6MGKjYbeZr7dPu0zYzG
4MiAGBPPvGkVf77KnauR8v3pxD3lVEjq9lwgh/UkJkoOhVCzYsAReNHxynVBtnu6nGHzgz4Peaqo
35VXrwnMgSHoPjiVjZEGaY4BS+Nf3UvJSClHSXmvCInoHtg67vy6aujwqrqDQvveZ0icCKqrELww
z221ibD73U5VhT2V3Aum+r2FPGsJT2EYKOMaUBUZiLCAuMSVuVN8VHrWKdKte6RkLYrVuEMZ4WMQ
VcC1I4/nxmGtlC2mHmaXghAVT488vjFoP8oxWLuCZVIvIEurF7OfYUFOkdwvRLKY6t3U0oT3teky
JiOSHICE1LFGv+0ZFFr/xzc2H1gITei/O9lnxiZH0ixrQofcV/hWRw9vdTteNcMV4leVFV/J05H4
amP01/sNtTQwiZgUzGC40raE2dyYfx8Mtx6BQUmviw7TTnk/vW8+oeTk76j2DOYDv15JbynsSte0
LJpTtU0zh+zikWmQXDAUiIN7h/ZMehJuozhDM+vLc0Uah0QGn9USg0Dui+Gg++jb/7UFzbBbfDcJ
bLpyfnDWBa/mzS4BgNNQdECMXBHQiOKAwdDX90hw7EnK1wm4/NDd1l/knKGGT3waIH/Y4TC3xUWX
25UZ4Q05DGqttAfRrtlyo54XHa1nONyw/SRNUs4h0+DrIw5bIDjJz0Qq42Db01BDlXFCZKozMl4f
pVwZt16JORXiXM2QHQeEuhpiUVx5Q8OOviCFzS2Nuht3pe6LnOKuzd1gOt2VFCKU3tOPRE25HoXy
L7W0yPkGPo/JT0Okk+blkcm8Dcm+ntI/n5mEy6OYu6vPvDjl6ybnRSA9MFr6+VimcvqnL6ccd95w
G/DAuJeGB1LBLKo2A1lSCHjkdw/bbLpZca6pbfl219TEf30olMKXY3KK9Usi8yTBzHkH+cXDdM4E
EkGAN4iMKW1IrUjsf15u85KA72RAletynK5u+RpJC0GRN0uT10CCt33ocsTGSjcue6DCx7gK6PiF
lBF1/q52vx9KxKdgw+vgbMdwYp0l4I+m3n3742gmDgS7bLBFPqE5pLRJkICiQni9G08HpwtSqWJU
jxLfe/0+jhQcf7iypt0lk19VDGUY7+MQ4122id1Pzzie80mrzJhc0uXbjXnrBCu6hPXlo7Aw0Qa7
A/CW/+1d1ReKhWj2CPoYyDtqvoVeCAn1u0YfJjFnWStyOOrCH16JTyoFpaSaA5jngVxbXEOXZDC5
mAZwefRUbSouwfMZzOR20b5bv5bFAfUIzcGcgnqd5v05roac/yy9nl2crFfXWFA2HWim7M2m46H/
aVuetginCrWfwt4vyg4L467OUplgKpxCtT2uDsOv/P8MK/k/bT2KyUqZfb+RInT+CDAL/Jg/Tid9
70w1+6qkwjJ2iF8fNVTlR1OIKsW+eNUMIy/dGBgauN7msKtaaJNHPjk/u5MuJxjWjx72Og6u6MH+
hlr1AaYspFE5I8+OjXhv6KQ3HZ709ZA1PSI3D/ieV/CCOvt/SnVECluG7DS58yD8HVwr5GAXus72
lLubGmAsARoAkYFDugcE/Y1hsjhAJBy6goysNKA+YjgasIBdFILaRfl9y9BMaqWRp/sW0FwvQo7E
L3As3yUZeEsvxVJTpZLoHpg5GciuCKRh6C4vZ36nEDBn/2GEbL57heq9xfgaQn0VOad58EK9lCeQ
EyiGiNgO5mmRON/DYRGqOGDwb5waY7yNo6OzYFZzV8jxfbbcCsXG5/iSjDBRm32sAkTvNHQcxnGn
BhIxKsIgGuEw0JnPrwhQh9DxYCKGECQiDZcAcZkXoKsI+rwTJPVcABkX1Q2qi0P68gYjBPMTWDKW
Qxghnzz/8yubO9sFwPyQtNaANpE4RDvWA8fH0kX3ZXge1MBJuWmnONY1zJZYeqLk4hh4oyrHwz2e
g/717pUTpu+5MIOk0krQNVxbATe+w2Cd66+CUuiwhF958iVH9Q/wli+PqnXwrgQ+9eTYqz0Eab9Y
Fa06ZVH6Q5MrnO+X6gXHH2SUqa+bJAdA7BR2+ltng/CgNg2znesPqUviIE+SSnLuLBaq+4scjfBV
SGZNEdBAFvUiFlWzbkvYQlAy3G21Upz7bSCRaxkAa5qT5z3G0OId6DWY3PAySyeBoGCHFoqRuHqw
jtMTx51l8ODTDtqJkgazL+sDYhMU8uOl7Xbnk/Ig3DZPqSr/P/rpwLcYB0kQBO3bxp7NbIEQjhF5
46Vb29/OvmDhWzBmYSyVQ73fSGYBIK8gMo2+4qjNIf5G7RZKTibRy/gBaBh7zWJxfaYoAvHThMjN
uFiI17H06AL4GgpiPpIXNGtl0iGnYkedPuGQCFe8z2Tz54gmdYfeUnkI9XYGuacFuzBxpLNcf429
8l7Lwd75jjrSAOhT7+M8es/a+DTf90o7WQYRGtQUxZPN1pm08vgueFpqyXAtVXAihyATSyBZCVhh
7yB8Ut4AvpIFnLF7YC9jCn0q2Ha5ApLzPd+fioUDJM5MUVKLlfqFufJoBbTR2ss2SD/RrzeB6dbq
j8aF0jaSNHGgTE5dRQL216Uxdo2ngZgjiDXekYFwKQYjaldx8ph9KlzU6JeTFSGjFk7sr/V7JHTA
1OR9UgcFMzUdNPa1JYm1x7rmRyznuOKGZ+DcusFmkqUgDqYPgjXutMcyuhyXvKgHykPGUzKYiBCv
7IkSVKtwrvfSbVvMHfit2I+Dw9HntrxwxBF77BbdIGsg4pxErIW4oFAGMADxCrQ3mBWvGYOZoCSQ
hQ4MCGmI+qe7uc5MQyhb7jZ5bPrPkMbcpAh/MuitZwlt8UcxUp0EjDxyinKE7BoSGtQUmi2zlnFk
nzvjSb2QXsElpYADQuddKynkSKGtaEF9N38c8/MfLQKz1OWDRc9yehNiL4kZksprA0+en7RDPM+D
kAU8BRKFc32RSmvj1W1KjRlEy6rClOTdmgOTeGC9EAPOr+cGY5Bbt0Me/gBRwYShtiKng5P2AzJl
6HPbWBGWR3az9vsd0r+KNQXo+3RMBDhh+GxAV1XwZ6rRk4aXexnP7VjvCkkiWApooji3txoTXbQp
twKputN0/0v0u2trFR64So1ZJ2UqTLmJlT1RLLC+znprAWwl1dE3UtfvLuoTJoER2hzBVmTdrHPW
gQcdb5KWlbpE8iersLvyYz5waXbz8F/h0tm+Xj5yRZ9oJDX/C6Gu47yamv0IHX1EUeU2cl4qjyb3
txrU8qF/ZQQB9pWxmkTpet4Z7RDiBLOp5F546VuOyX37saVEMYT1YT0Gbfp/0me9n/JcXbMQQSar
opuQJc+hLMyBmoSHSAqUJSWZWhR5cU9391uMXvZ19GtIAwdZBdolaHDOTCFKHVLQ88IiBXIiC21z
t7AG7b5AMgur8zx9dmu3NDpphXXRLjc4nwGlTGKqFGT0l2IsmwW2lSqac7COML7nth0msZ6ZJwfb
TmTJBfHQ9E2WkhiokVqwlSBptK28j1cJ//253972XJm2+M0N0B7bRnaHeZdk+F5tw9fnIriRHigH
+8PJODyiPOTVmHlpJwwPpbVhTs9cnBwQ6hgNZR6qDYGNKWrkpCGS/K7uQzJItIuJY9tQ6GHQfUJS
cFtezT1P3k4W7r8Q4f+7YIjkN1cRjqbOrtrqISH9s9sS1HaKqBAMuGPQAqy6zkeGg0etniY1UInJ
2eYS/7vMMz89CpG3ZH+YXB8kaleFGC88ovvmPLO6ZzB7z79Hm1SzImsdKd5UMds2iRKvP+Te6eaZ
EsGzdoWopYje3Nj8+jqAtM9NU/bsntilFzenC42g6oo4/zqn5ytid8hU2IZccv3HJ0nHtbnS4vdh
53Tspig+joycFqMk9NtZkFOm7ly+EAK+GWw7FoFWfX0bHepnOVgCds4DdnL/bXJ6FzrB803zSvnN
v2n6mIxiSE2OnVremiL3uegVLG0pRWYOkYjmlKOaa9loWxBzogZOTIvn2OxkIZKZg8ANWUHPxA2w
18eRGZcSIsyPJUhYInMPGkXD7M268fB3xxoq72yJo4MS8YptBaVLog32bJOVTupQCOJurtuJXlHV
H7BIkl/wpHxF1r6qnXHQjkqmhsobm2lNn6v/RePYNMgn7Je0uduyse18j9+/M5s7/9mOX66uchO0
hYxH5k5Ucnlmg/pprCivTzCyxPu5R6GrVdCzJrySfJwrG+BPBO+dCwPLmEAduXm5eEPfhXhFbHKG
F8efFOJUPnxzbfHC3b4S9wBGRXSV9fPBUhrve1b5be+4ujQ+O0eD/EAZ5M8QrlMMypHSsxAkySMI
GWUe1VtOs7JJ6c8xKhgi6kU+2i62DwD89nGtFCYJoCmELCp4YqUJoJPMKdgUpZKd0WjfM+lN90yt
OLmSA6ota8ro46nv9PbRiKxl5eHmwXMdx1j5QPKuv1angGuti8t+94vXz77STLnfiCzZzq7G6qp2
2QzQVRHapylOEOzKeDrTPZxBPiPqc+4TlcyR72l7cc5w76ROCKEm7IyIW9Io7ZX6euC4lLx/1NiD
IMh1a7BMUHhwVFbyD/eYfOhN1Y4LE4rZUfjLbMkellwpSLxcW0+RqMuJFGZQ4Zwm+PPtZJxmS46J
mWM9mjmWPtH2jDDyiN1M1M387pHUWS0CNZwHhUxc3iZu1c0KkWAj/4ETp0jqu+mTrmYfxvzYm+tF
1+y8E0EwhYvj5QUsZJEgkmz+xh5YD8MRbpr2qec1QHKtUteVgrCoXXzZfV9eXKwjZNC1kYtXCdbG
yJoBC5y62y0WRxpdEM1tb72TBRx8i8sZXM7T8Wtdb9uPgpo6Fpv7IUeiaKDhoy5j/skHL8lM+nKG
z3kaxXFVSA7b2hnc5HRot6Hm6GJ1Z8kwHK4RkWpZS5quuhC57lxkCJra/3ocY+wSSDrnRjYMl31u
1Lf1ot8HJ4tVqVfB/HBF+8qkDvszJl8mdCwD+BUMPGEybNmjabr23Uf+MYvW0pLdvh5OlmUp0Q5X
AKu7gqJrL/8iPJb+VTLFnK2GqumDDhmdXVhSEp78xKIEjvMHVmxBw2Z+ijrVgysrEWoA9aLt5Ahv
ouv5X4rdn3C2nmrRZ0lNQHz7JYqlRvLahxkoTVCyJvM2xv/AxZ+K6iXuXaBKC2fPEaFm48j/ffrY
Lemktj9AlZJAfLENH3iFMbkfv48Tc/3OSrd6E8eSLET7zqij+w8qKrI+7So+b8K95m3H+GzfohCY
zXTkxzVLN4eKSKAUrMU1pcT8DRbGCBs6Q9SEduKBrU7O4y2XRx8PKdqs+h6ZF4ba1PmMflzMpme1
pvdzlGtfRX0KEjW1PgoHU8rkBTQ++Ka3wILKktL8b8v3wrjitszS/dRqpC6XWmbkKPXPYyUBVkwM
SCQdxif+ajMYT+7X3Q2b3b4Jg4P4LZ+vKG8CAydMgQ9FsshzN/pmYK8Ek0lJ60MvCkqFLLxzp0YS
welxfAZxXQdiwJFpgS6snEKMpsc2QPqEGfSvopa3W7iK6wd09bHmD12YKI4t9ENErEr9QmCcv5my
7OLf0NeXkCqo3Tl8RQBARSzyWkh8HWqPAOUrl35MUmziQm/a12UicWjQvKdkrQ6yPEg63VWUqQSV
BGJ04T/dQtMxdnalcTSNGlILmwzakvaC22p5gaFqdSZKw5gasPr8gDrltbyymFzx6cR18HwHFjk9
2uWJ9Ar1Qu1HKiF+8xpjkWEs+VqBsTHedYGAz4VmSwXAdUHw6d43Xvxx5b4ZfyRjEoSeJqgW5QhE
Zik3trNkEAZGtNpux/KhEaOSSk2uEuswsmM76BFu2pzlvZ4VFnvg/SXvaKnmd1PwMHaCRi1UmaEA
j2oBOt0TmkR2bIVZGtoyZobKs66TXkc4i7jF722chvFjR6pimCB1bvzcXA/vRaBTTe7ChvU4bGDl
xocC32NQ3k0fniw29p7Q5E3BhuudTns/tpclMjODZK8jgj80GzZLMrrXBtUTgaBIReA8Qj/aJKva
BBPQ1p08XnlCwhKDgiNIEe3R9gbQ5l4UT01KClLqcjSA574KjtHcfgf2+dAI9dTnvp9msQNs/RMG
CYkBF+QFh711hmE1uNnJvHhuJ1YXVp+Lf6UT9o/osR9UEBUXTMaU/s/MGxRsO2ra0RHcqEZ1zqCp
WZ9NCZrXEd16KO8EpAekXW8JXfoyeXLS6VHP/naTmOnueubQxDM0Vr6HZcQZTRnD0Jg8RC9HH/0R
KabOJr8UZEDOTH6DnOOSy6xPwJ0swy4XjauOgz9dmCMN6RDcpbbeXqIwGTuRemLwM1yeoTHD9gsQ
TYXtqBm9asYz2ckH+6SdBkvsMclYsIMjAMFBHxt2gszCiJB+7NRoPLa6SuZNttsGEpUKWk4Emtbk
EXpDzhbFbO9JmHw7OstcIJR0Zo5F6F7TXPkOJSmh4TWJAA0d+HBvyi7n9F0lq3aYCNk3Wip3a0hK
Jijp+98xykSzNv0fGh0UE8Lm1dhSYXaPAQaYKHLYSKPaawGnNGFmuvC6I/QShfNi2AktZWJh89CD
DESO3IfzSPMSlJrQ1KgiWf4NC506Bm3cNAffQREbif08Ew7h3gQIyllq4LRVvkQivMockuM8k6mK
w8jicggYOXeNkh6AwqHJBTIb9GiPk6KLP4IJBKUjW0QaReibrq6mumFJQwgwLfHCz2NP6COJPuJf
zgK3yMEOQMVi17E+BSq3sYjK1fAqH6L5WQtEUVhdMNI9SCbAWPAb+dWkn7nC3POXICS2jpJj84GL
YgzU0USGCCkWn5AkOP3Z/ZiTfUbBxPDkaLBgX6T/NcjODGd3UoB4KPjPFeSzWqxdYPHHwkMrJP8v
CAPhKfzOscF6k/q/Frxly7bHpjd6O5sXqq3nIzEqySIBMJ9dbkpPatHiKF+y563Xg4jHCSzgWQrI
3n8bCcMjlFbnePT0kbQll41mtysDLhMynRY7cN3VLaeZatopGVep3MmVkR/tF6rd7Y8hCgjWhK3X
t++uksfkbSQyXR9AN97IJTxAcu11ElZax9a6/dsUoF/VGG+j/fZdCchXwTTrApMRAZ1GVLN93b85
JuO6lA3HEgHnt0Z3Pqxh1Rbv69nDEy2tEvfKKpFfrWghoDamFDlZouPO/UsAZAT/ZTMwGGfKwCvX
COGYqiNS+rKoUGcmDO0NEN8540r8k9vfgt8TFzBN3HFfStSf+7J5sc1z/BfL24vEEDOC2t+qtrzQ
oeS1EMA1NUcVg7QJ5TBJk7U0IBzACM673UyopEUF/0FpXsNPZJVh90Y6+Xa2WRc1Qd5vNLCSFaJ5
6rn+AuJh5/leXCmVfaAA9gizRnpH/VpWhpkAMLv8+RnwRdmN7JWbq6y/X37j/eIoBAnEO7chaBeP
4i8dLf7t4CdlVc5xY2gfmSESI6AwXZ/YWRwiPkQEnyuEdHhGzm8IfRyKANvbs6lxigcoB+AXK0Wj
eNQnUvZgH1ALAK5CKLUWnB4NvyLLHri4T8bBW09oP00PHg8tOcAD99DmgbADOfIqc7fFTVUMZk6g
a+P11OLGbWdv+nBGuOD7uHn1P/Gy6U5fT4O7ZXm0RIpFd4AOfj7OmXGn+BYCBCpetL6i0deEtkuQ
6uvRHUGVtlb4Mvrl4bYk6XsqscvEdPbtt8U3ulgKPyV1E+tmw6MAtToO5/K6oFSEtO7M9VhaN3Nd
fiuAJfhio+nG8HuwuEbnbQq2gYzl+JPWpyOsmYtbfgSzwSIL+mXLpNOnNDj+GBzj1JddE/RcbSa6
v5xWglQ+sa1WGywX7VehTKL45HhaJTb9+KC7V46wij5V+3zr+bTOxrbWGiK0K1ny4HQSlKqd+RKv
JM+JcTwgubZWV/ry9mGbqJOJ4qrnbcODX3IHWSpTyD1flTx1AauIenRvkQpC4ckbcbqojrcFvXHy
vT+1rQyLR8qaiG8ZCdpypwNW23tWBHc1tmPBh4Cj/EBfWST08vN1ZEMKYWOWdRqlekdbv9aae3V0
pRu35/GW6RvGIZMzHrhqxj+haqQARcPWk8CIsHkdLx1Xa0S/ic31e9FVYpFr8K4WekBt1sBGRXWR
66kVaFBr1btIkKCirngDbd6xLH5cQMh4s57dge6UTfht4UOHS1N1ym7cEdc/tA6XUiMtnv2GrdQE
O0AbChW0+uUkduXgch5Hu3lC0/Tq8852XdhptWAZK4VaCTVHN4QAhp8xnlcwRuasuU89lQfdNazX
WVcCDX0+ZHlpQ4171g7FQfqyg5Ky0XPcG48i0dxVO3b+vVPHr/wev+g0C57U6hNYmryWtTWnuZr6
4gJ/o2w4gwRBwSuUH2mg0pjnJSN2zsq9FNkzhdTKfSc5pzoIp7v3im406g8asaQOhjH1Yo6ZqWVr
mbLOecefKyIRRztMINwemZyOMGK6w2HhItcnUWXofQGUmx72xfHnwI67CqV3jRvz3PBia4UriN62
dL597k7KoMmHD7bkJRzgWvTUOMCxXEekKoDFV8bPJFVl124Y/9HtZusUvkqkV5K4Bvi+OSfyNCI9
nfZZTtoOmGwEH07dz/tz4Lh6ZqDfCRVnWVaZHLsdE0AqTNVJJZhHcUKXnha1U3PUBZ7K9hTDIQY0
c2UoxKGqGEmzOlXAF6iV5x2wh0mW6UrSt2p/JlQJ4y/1SwRH2YLknfgLwzFTA3bAg6LQ2H7hzPdl
9z+kF5zES8deiuE2Om6fMqgWHlw9/E43aiZ4kCap7CFD0KU/8PTni483UjsZF8Ts9gngMz1nElp3
fFf5uiRJNOsVM8/cYjxoBxd3dGwFh8gjRGj4PTRMY+FZRj9+qfs3odRvEQKF2x1g+PsKZhqIy57t
43+Pi/GH22pXNghKa2kLl/LonamdaEQKb/QanZ/u6Iw5lVuayLnMe6leeS2JsNDBSR5G5yIBI1Fm
GsQ9Y3/kEhK5kRL24JF7SYaRBamyb4BkvwjQob51GjOWuQ6XLzPCh440ypXTDTg8DBgNtluL+Zta
E20v7dH5Un1BMGjPh4XeyNJOZWYD+N4oTQ8BbJiJux6TL88TdlXSk4b+dbqUPKo8qfylFJ2UVcct
TJm6/t/PYf0sHX1v9rIwd0k+QUlS/OMvK0KEBz0giEa2Rgwz8zSr9ivVD00qRiT1Ch+FWbjkKJta
h7YVnUzuUAe5BM5MbHT4Lx3bP1JPvnYqrRKe5aQp6yRdKjOiFwWQVMXTgdDIoLBUUrF6lUlcD4Me
C1wID3Pj2j9gA1XE1Q/CASPWPN3qFql0hW+0Musu5gCx4fEGLargRQ0IentRfnMopvST9H46XyaH
zcR2KfTCcwYIeNDvo9ITkQVxN2B2vRUNORPLeJmaorSzCpKRZ0XN0mxadxL1ebEdorSKOpxRPh+S
4nbB/IAxJ9EosuqYRr7rK8hzRBm3nhDfjlLVEd2M8cCesep3bABivNnbixtLZKcnCbWY5Z4rOtJd
PgZgkDIyM+ZinKw5+3ndnaiiLgsqph/KK8GiJxuTVUoFKj5kUTteDXLJwgaHPqGQZE8YOyZb2wNc
mfZq/ncUh+qGXQJv6Cym+6dw7+2JQ2nVDW8EQz44JSAXnIp3qWrXK+15hItBMJvbwMvqe6cjfWII
cHZmNKtp1LNaCBt/aLZeWMTqSvpBCco/s8ipnow9RCgXWcPTHs/vy1/fOgVwiCwWP0O+jxZ88lew
ScJPIXknKJHcY2tBdHIXVB6qLQWS0oFWUHQ5tWcHVwdcsrA+hf1KQOzCY5cKC4oE/uJqhpRW7ls6
mAt5dM0Z7yrijUM8WkeR3h97jUlugsr3QmWQSfwu29sxHQMsBEz5sAqWOfZHNQgJCHj5xRqderyD
Grs/d4cHHV4Mo1AS/qRy5BZjeQ15DI4oLVDN1jc1yVhaDJozwiqtYjha75WfJuan33mVU2zb/EwZ
xurQsAiBk/KXdrJFbE51uBHUM1yBIlJ4BZqmRJlXovwf7EcFYcCxsSlgbbgr3UJ0nOBgzMr8elQl
vKWR+OqfIEKhY4dHZBLsBbkxwfdLYdKgwjVmTwE3oAi2iuMRoWTGvr2IuAR2SCQ2UkyBuAXNE6CL
Mp9MSu29iuFCSevh0E0toTVwrmNDheA9+DwDsX4EvqV5Eik2etOPsLkhw6MaxhDp5yxAWnZZeaRg
kXOXJcQsAoPn1EIlc6AfsDexubZ0sz7Ag/459i13qjjfobfpRGnZks8KRGFwAQXW4rxIqFYftgbu
rUSGNz+qzVwSfJZPHDjqvFoLCq4QCQJxOEx6iOFuBmWapELgU5H4Jlyz5nqVHLG3bme607hKMKNL
MggJKPrwm2vJ/O3v4cyhyEmXV5aGDhsuncKnvsar2ztjJutwG//z2AZ4DU8czrSMPR/wDl/+9Ll8
Qb9Jhm4YFncq4r4viij2qNKRdBkDid3R+e3hNqmQYPJYxG0vticbIMm+kUSlJ2omqmjsXSQV3q9P
qixN1J+Mqooc8aCE6EXtzfApIva1ZNEnb+g5PvJQqlIHJhB+cn/ljdl+uqcG2G1QUoJWKYM5oF/7
sWVGlJ5QDb1IlMpRp9yn05oFMOZibjbyEDg2Ck9rO4LOcLdmZg76eOF4Y8nSvt3+aFEBsM4kNspM
dCrB7ZEBjSoD5HEegPGXy5BwQqdxPEBBhtQeltx2coJp60TfgoQNTFm6UXLu9INU8SfjxaZMxvr2
Qd37CWKsVxKaNjuiF0OIFeaUong4BVq1+thn3Lg88S7ZcYCXnqQSGsPpd2lIXpSPK/ko7sCaOfU0
9d54h54wvHYEBn+MhCeX34XEluZALZv5Nss0G3gV12mEJEy81Xk653HIdRjRDCX67jTtP/xZSGHb
IXOA2lsoKS2QuRztRD9zNXS0E6QR6ldqK4ND3M9Z/V8WIt1khTwyDIXoOc7/19u9Vr/3V2m2Gom2
RdPqxFbcb14SyOdEBMUJjRTBwF0OVGe5rIdRctLJKqlIvZfI1jACBlOn3B2KvwQAPvHhahnYwUrg
70wy8kOvzVCtuUvV+xeb/eLi3CGARWwpZHA26WYIxyjpbm5c9GJPtsUbjhUekFWqerJRqxGcrUev
wCTdn28XjqcN7vYVEgg5C92bQ0yhNgvA+c62Y5QSxZbEOcUsvwaYNH+8ONSmqFE9YcWot/THoo/k
13EzBPZcgZdzpvQ56qYV9KIYM5f5fRGrrRkYAb8yQ6u8DTZZUkvPaUX/bSkR65meG0urqn1TxGEg
AHR6GX9tCt7HGF9EUqE7zwi22tIZBtvP0dz8jfNIsxIiVoVvLWLIgsVEQF6uD6QJ9H6D0L4cPxQP
LQzl9SgfJJfCZmNyvf1/RnAkexj294tAezwL7K3R+EE42GQvBUkb24nNsA6MKvoJof1sB4cVg8Hf
W9QZDkVnYhVMMpsR8s5FoKc4nh8i/ghvoZhB3ed8Hlbzp5p9qqycR2t67owMT8B9pvnDkTjaGQhs
nf43/of03NnbY8WrdPgHRPPmf/78xyq+8b+UJ3zjBsck46esBcKi89OnLEc2Y0nPWTfrk24f6QKh
doNfYgDh7a8+80neRCNer2D84cP5SPJZEdl0thncksRvqjO2D2R0YPLkoN2wzzHTSqbVI04Bw3Ym
rSsuXmQ9nenlns8neP1C8HSh/4i0de5bV8nyfIdDaenp6XLP1OSkjUiWfqAx0x28FNCfoZg6N/T2
D3qM7rKyJotrH7WWE8pMBxwvkshJm0Uljbo8NCPr6fm+VunTq16yLrS9/XdqH8dLRG19t/l5sOmE
MExpzs5wwMurS08MpHlMsPY2Gg9guaZ8LK6A/vQOu7BV4LjGAhEKHO7uVIEt0kS/ap+F8MMwT6Au
6eIrnpj9Zc4EkB9IDDtkhB3N8d1WthWrqxiEhJwrwkR93pozHzit5NQ6xNW2yfWUrrYLrkjc1P6y
aILyEKyPAIChoIucDoLxvYJ/BuNcg9Kg22d0EULH/1W2jkWkjq7MTyab/KfVQ2yJwNkyasKHhf4A
88x8+FgOxO1B6xenIOyRQKctSTCe7OKhhRokLBxSgs6CyzOPgReC+H1MVxm5HanPojYmRv5kv+Ws
jiQc0R/WGthTteyLyUZdrpZCVkte1aaUH8vAl0r3VfDmwS7Vfgo4m8FX3MJgTdEifgsECb2CfKY6
hYgzQUiENTvB03nvvSvR1TAHwJBU95zEGyOnhLEjuQoj05W7SSPInznEs5jZJ2aQY8tNdrIpL179
U02q0EwYF4G6DP7C6ENUOfDaIKlr3Wj/eS1cj0jP+gHfAF2LZmfS0gOqwTaV2QquCq6qT7jK/g4y
2n17D06CZqIeqfbt0suEbdA2hsSE+8loIYjIWjtTCrcovCTQRPsry/IQihaVQEKdYUFf4PiH0vT6
07nSvIS47dHEQSlS7fOUaYvmD1bJwy9A24R3pz9wx2N3oM7z0seqw+sy9y5Z6xYQHmwjVVA3AtBm
xyWaFVWwG6sYt9Kir2RRiEGlv+QX3arbWUTZNpX/ux6bQ2f+/KqVI0/E6fa7jHZeJU7m8Kebrweh
CjUflzoNlpsPFUldhOxcIOm4SHLgmOS3K0pEg5nGVIXcgTQO9VudQE4M+H8Be1zkYGlCLtIFZgQX
rdlCjDb5yJRJ72s9OPUVU0J6N4SMONCWo6T5F52kz3Q1qdrdfzqROs+coo0juqWafsOjvRbvmp61
c4x/5/3AfNOL3WYbQeImjQx/R1FnM1ChsJsJQpt8UuMrhRw7N+NXr1Yuvo/xRPgj6YZer3B3Tqjs
9U6O957JiqBMcjxWPrLtTqFRWO4BFav0bf8t8J3PMrfr1itKs4GnHTLdWtXBOOVjLThD2w4UqHYi
ZpZZQH+HFb3jAWTGY2vRQOKonE9rAlRuR5NGgw9zG7RhcOwCZpAyLIiYv8P8VAkWf+K2xXA61p/t
VJHlxQzNDqbf8cleXMgJ1DQTrSQvcKw5WDPSkOhLDhIdVYyoK76grdwT7GGKGiDGMXcNuE7fptLx
IfHNNyVtq07I99l48HVKWcIkEIjW7MiXxk5A3JrqYh2WIJyedkTmkmcpty7IAigrpbF/v9+fsh5Y
tzm+pT25iPa5kQqDKLwyFDNfiKOaeSnzPB7V03Nu7Ks+CBaqmJDaAPaGZ/CYyMx7sacVCYODDnuA
6rCxiM3wSBT0ZeHObqkRByWt1DAsnJgL1zzwwlZhH8oglXhcoxLBpemQSg6Z+FCQ2BAv/uuQ85nF
55VpVUxvaLhBV2zx/AaRzo+dg+ET8ylMWRBJMlhvD8H9EOSkLnNOg4ziqpka6pzEYIW7RcYqD4YZ
9qaQooqjSIJRxzjgf9TYA+mwRWsEu2E5p6jrTj5/8kAVqlnILRdVULkQtYC1uHzgaKFs32JaQIhE
xm1woNwBwtEMtC0ES1crq/FWVAppzRKi6DCJqHOoDSs1h0DXW2gFvdXYY/di4RDLBa9gCrAW6yEd
bSpSV9whGSojMr7rmlZdKKtpfBtWmfoHGglfyvygP9YZMjJG06ddpVfGTLxd+ugbLy69jHklpA+A
xLB2RDzdzlT7Ajch93kF/etiZT9bdsDRjds+Ll98HLhC7hCn+JJwAyBGNrkOhV4R7PYnUYGRC1ay
xOhVOo4v7jnMd5NJe9uOZFzRdT/99tGytM5q5zLZSmpZKdOaBe7aIRjfMtjicZbHmWcYy9D0RKB4
M8CTNdH8OnTwQB8vfwaHQMBMs2A42uaSmeq+/hviGzALO7vDitUE3OH5p9o/iBPABsnXPOtgibM4
6mXlyoce1Tsy5LqRzJuXik7pPGqTmlfNBDaOCRThV4Aa1fb915qVoLVVUtNbvmfQwMgUTq2NDawx
zze2WIHIFvkhOW90lOJ3We5KD3C5NRnslAG/uKPaVDTCeFHNrYdAXbPD48T8vfOZ9Y5Juno5Yl+1
hikgUBnAO4I6A2fsivhNCIuKb6Atjf1M+19lwbvSlLFB9Enwem/vD6HbImSO1Iq4WMK2z0j19vwU
ce4xT6dJXfjB2Mtfo3FIa3r0xqlXx9HNDX2AhHuOoLFrbYPIDLEI1V+k/56uA0SKa+Nnoc4JW91P
DAib918ay0HnIaLlUr21rPpR2YR6LBvuHcFRplX4hx4SKL8C5thvfhslGOFmVnmQkeOpOQ6AUE+I
A21gp0QLMJ+4186wFWCUigV9EShipeW5mHD1svThvpjrv+IJp1ptjxEC5WDNnvgvkxIX7P0tNvSC
PvjZX+c71g0C7lae+gB48Yu8lKQcoSnmSeaJEGUiYO4Bg3lbqYdU9bDBKy0sxj3xFiKgBrGh+unh
3/CpVdVG1YPxKOcDMTRYg8C1QH+2LQaNJmbDLUMPyWlewNcjTXPThUZaqs51lI1aW/cu5aIR8xfv
6c3frx0f6eRNC3rlXRUwSVlr5Ep/scXNKVTBnL6YRmvBiM8hG9PDup3XPzKC2LEtBm2rwYm4ul/o
zfWz6j8bA8YO01ycc2q8H9QlMmGpMzMRclU/SOAw3J+7FF1f/uY9o5ufg80jIlp60gVFw2d/5ZUs
r7XAbxZ3rN6fKgb6G0oE686xoiWWVYJAnMYHF3nD2oJmPbCyGTKjkPOx1cCMUsv+zRxg1mlwD4Sf
OvfqtHmSbnj6UtpwBSX3FplBVAhYi+A5eOVdXHGEzGtGZpyG9IwYmVS/1QlcHQ9IvOcoCnEvP6VV
Y8k36H3oPrua3wct1OoSJ4+oTFmqBdOtcq014eiHCAWGXZU01IOX6CxEYjL2rq7KTKg8jdlEQzvJ
QJdYST8ScIzohVSDbXnxbL2mHqEENMnqyc+xZxzhPopzBL/zpTHhw/cb2Em/+5/OYDDpHDeE/Jsu
icatxwC15rXXY/HpH9L4d//1pL3+B2OuyLCK/A24GJyC9OxF5E1e50G9IB/kSb9mCVXqxSjfiEhv
JmltPgXJ5BX5GQMnR2R/Yx1dNIZ8OAQoP28LpS0tRZv7CwYj+YnD0sVZ/BgYdRsnImtPfnIdJRKe
gRER3YZzjQDnoU9PWZigpIYDKeC9XL8tWJoSU2T+7122bM1M0Jm35DpV4ZfX5VSEk23wF0McbY4Q
W7CWIayaNMlmdb2z5YjEll2v+V8mE3G3FC2QYjmwNoUC6j5QXKFxf8I8vPYIKbE/HTT+ztHNj41h
7NY65bAzg02Ox/xzaKz71ps4q41QNK6eZaIrnu79/MYvtRdccTaizQZo0eCQtd3nRBivgusq5iTA
PTy2Ul9uopMY7glciB5jD9N9kkolCqP5HY2EkYMEAsbtgbo8evnVzlRJDxWiTqOUrAg/2jRDebIo
8T+BeusQcU675MgZztkYmGoe3C49a/Y85f1CZ49HK6i4Xe7F+kQsbqwZwypy6zi7H8fSc4hi/xi7
OmDbvTxvN2W43cEKbtI5nnBF29in+3j7z0xPOrtQZPOv4ZAoLj6K0LTOdr5e+IWUXhLatNW0erhc
lwCTcAGndFHcKDG6wOAl/xJTH7yhVJ1R7GZNsiwynspewmIjp9FEvQsPWztRYZ4kGixwZG4AFwaf
+i0AbBtIKPRw6B9hRqqyfTvtgPxs2ajvbS9nskgOR7Sy8rAh/74y6F3LcCafYveHTnBPkTyBg2k6
rYQiBxj5DRfsdrXmVxo5iXuofCnf9Qro9i/Ho1SJk5luFYxMe/CSNG5Mm7XdWoXviFvfJZTJ9aEd
7PC8Ap3UzCIwSPw+xnerK5F2TCSF9VDu8GC5/rQXvLwZUgDXFpeSVbJ5TXu13Zy2l/gABTzZGcEq
Tr/QkcIrEfe0KyFiKbiT3zIh1Jak2aY7iSIdmQ90oPAZBQ0YuHRnl44kL+BUejAILr4jdEGwlNec
MF44bM3WoPSw2HuK/dEfPF8jGnb5cXiiAQvD/NOQnhFTR+87wMxZM4VqE6TNQUuZo4MnGzeDtBy+
zAflesWHD8gSViAY0NUoJBKRX7494dtnlkI6nrEWHAHcgFC7kf/WSmed7Hdq2+FMcB40Q2Wy6RZ4
CP3YYrfuBsX4KqB1iEY/F3yDcCGn4m6j32zbqD8JAuTAXSTsJhI4pUNGt9u6Mv2yXqZNEfDXqFrn
0EP7mw+z1PrL9OuDimEXto/DiNagVa1vM1arkjikYLxv2UzAlcuX1gRdIdzgjN29Zd08Ey8wjJEM
1d3z6vFeFg0f7KVPwBJDi1rqxo3nCyYsxfcpZOcascNVBnV1fV8SaE8fz/b6aLWt32JtQDbprlC7
xcOI/HxhfZl4kFrnWHayZUdCLSJ7GWjJXeydf9L0Sks+L8yRbmwH2P9pVO7k5RI1iRp0HJNtMgrD
qAMOXZm7XS21T8II8sKtA4xrSKbK6qZHjclDqKsdk28vt+NDpfjrEVBUM7jaKubiBmjahd2ungOy
QSPtMljt0PDtENkY6uPO3gTXT4R3P8VQhREnYgij5lkCbG4Mdx4mZa0hCGiKLKpHnsrreg+YX7yP
g/CPl1RqdZ4eVvFCge4vMv2yn9Hl7wwGmtOxNdo+t4+xbqzklCo05k7y7VV+dUNtV0ykMnyJgss4
FwTc23KfRn6kJsklZnr+fc7hAsUTInnGy20ToGDwd6y2X7W4yPmOeT7UHCZLmp0dIWQNg/LfmmQQ
N8rYYpmk+aiuyfTcDeEmHSPEh5OQXI+CAesXwoGgSCUvr87sYYnkNhd44vX1wVVR5Vh7GQOz7Nxa
fWxYm7TledL5LnoWrllb5mT746ND33fQ2m4y2JmUfxrxTG6UsXjuphpcAsfdEn9ZacPrUla5+0Ez
Y5gWiIQ3kDe74yzMQx3ca0b4VeEpsK2kiNbjtc0XoDXE6uAHdo9TziRZT4LSA49sQeKZ5bhbnCtv
ye62cvJnV89eRZekRzbkqn9Zj0WSs46TqiTTsUtRzhYdfcoSzIHQUA+JSh5PKzJHCwmBhrrIK4xv
miLIoX4WCen5lPuIK5jVRbTw5XpPzqX7YS8eetUtgncnP7/uSmvRE1Psj7b7pq+6c52+5zim5wjq
7hd+EBq/hI0r5xtQhtprqhG1YVe5cwmkDPKQjEKR9EHbDV5kLsTq06ybpK55FOshl5+tJI0X6vXX
pXmF/fo5lWn83oABXr7HLXY9SZSyzxtIRLahAS+DsxgCsoqvc2ZkEatcZ96sJD5WgrXYcOK9tROr
RvNhonuc3WMgZfZNsNRpwHD/eFs3E2uvOU243VqK5fYxBi9POnSchJQSvedJ9r7n1DDRsOhMZnE7
zCq+2nONGxTNYf2yMc0BrOy502L31blpFSdPHf4APORrD4jN0cvZtdNSNlYOVLAT5e4VRevnF9z0
cZ/dDDkSPsRcCbKKmziFKk9r5q38NOa0383HG8aBXncOo5jhap/S1S6d1UVhyibf3y336PpKL5a7
WjLm2JI7HnhPhazA1AVfE5pPaxVmRPbtMb5r76h4HylUPgjnhVzrdYj7Bs/a4SaiFWRSWCo1eVC6
7sD1A0H4SNPOGut21NsrEF0Jrm11oifXontx11B+rB3Ot8o0oRcF+E7lY3hideUusmKNUstB4HaD
v/bClQAlv82yDvVnT8UxQlqWLGSSp9x82sDxok10Rfs9RLtcEkpAc/ZHVqpqM+BSzB83ysnuP+FW
uNgDYWzZ9MIWk3Bdh0U4PxdvlgR8gL/d1xI/oP6dH1uRvGjOx3EOPZ11/eDNXhcq+aM5hXI9GiXZ
aKEhsPKtFPmDXmoSNfukdX9I+PoH6GZGq3iuvPw8W/uVbd3YG+Lc7ou/45ovpQFapcBOJFUQNuVK
RV/5RRTncElnOaRgqC4HVVhCLh+fn80Qita/0ETyq3p5ibhWiOJ4xHd3YmI07PzLkAPUOIYEWFyZ
zpeF4jobIdUNxTiXAJDzgBhbxVtMUnj7XZezsnAMt2B2r3LVK/pJex0iSRjvHqPwhEWGv221tf4R
IB+3ssEpDS2fHXtmEgZO2I3ls9HjOoS5hf4LmodDSvgu/SecsF1MPZm9Nlm2r13J4ocvrxbxOVeC
ME6Cwo8bB4rScyPAz3sG81BkaZ1GJz1vMcIQaSWam51hk7XXkYFN1jFul59V9k4P5Kea1KJ5rNy7
0R+m7Q6K3W2cMXvw9gll1M70crZmx1tvKrzF23LHj2EjAzfNb506RKC977mCJl+7tGdmYu0i1UCa
vdEsdhebqLVq76L9YLY9ru/gQBN1uFL6H229zis51DIm7EB/Q7UfMrm/kxdcnxrK0Xx1l1XQupaI
jJabSmI3GoNVdA0pzXayezPGv4BRhFvM1CRsGZBBTTIiugBN0EQsFTNEjljoru7tZZntinY7/hcU
wk2cCbCH8wN3I6sr2PbIgq+ShFRjCxyPg3E1YVb4RdSfchUkdfLrV2DAz1E8jnJtwyOtTHhgRfBF
oim6kXyo36QMj4kVHaNYhredYQXXbkIOgv0O5BTO7q+mAZr0R3e9sZq1pKY5HfKZZvQsHpBin4xL
+8E/BH7QdcM1bF4Q0sBPcI3Dy+jZD7l244C32f9GWdL+cJiII41iscInOvldxEwstflqEUTijHpw
yPCbJPbytCvtj96Yc7icOKMYlTFY+Kjn44DcQ+w70VQQfxoGWEF+KWDvgDAJKSnYtJ2mQvDRo1up
ltRlYFN9s2Jlf3Z4J0iSir3VgJPKAUQgx/MsWz3zwsvuhmBtj1BYWfKSY9k4e7HMkGsuftwiDcWz
m2/pnUXJnzUsqDE1vLx9H5IUJzioPDix6ybN8Qe3meK6m0QpkAV/T+xIw9ZXcJRlKyTpE+B7Bbh7
Di5sY9hkXmAKjwmGE4+YmTR8raZ4fMkzs/zIDqCB/xOzDIt5zWRK5kXADjOcxjSRCayXYErt/MB3
h0wtAjCyTCm/NbzrE14/ry0z0y9zwr8PgS9GJQyS42mkg5n2sYorwhYVJ+o4/MXvzUmc2yTm7TJP
o/Nustrf0IFNAmjD4oMQqYdnS/lgYuhgjgfAoN3zMvqWApOMvMod56alDdaABoXa1oi1Jen5x/6B
QrqIY8S/AgEp3ozWCZXUYQVsFUCF/bv3i+e7jGmBixl3FZclTsKnS0MecD1DEgTbfq4KBJrsZijU
v19WOCttc06iW+ZxoBqgKqco4/VEYEgXgm7L/zdcrI+OUcWxfIBqV4DdtKjpu+j0uof2u055WixW
GW6Kz+T87ZI7DQHs7lnMXc0FAFli2tqplfYAOTWzzjPZWxo4mkzn84Y83Xo86YxQJ2Mn0tykYz/v
oKOqZJnRKu5ji6quXTZwMeFatNmdy2fqxKitLvEHfFSZPnF+ulxlgZ2ZXUGA9i4ovq4THPmwWL5k
XAf2+izTrucyv9ySOBcCJIPyz7666ukmCfnWQOlGm1kJ3E6e4h5/KwHGk7ZUgMZXzGfHZqxV2iyy
AmzRZm4+WN3Qc89/1GsASAvmdhvqhYLMID8wNiJLACUGG+prUjmwHrE/BwOTgYmEfsrlJKYLcCIA
448Q2FFaO+Lmwgp4MD9jRe5Ji/CBnWaM2SHdlVzkHzt7X2chvf9Xrsk4ymSF/8KHgAIrBxDz9p/M
dAeyIVWRN4B2N+ykmZBwpp0Iue7BjQ+cmg7iIXvUEa88AQh47gtwMoc1N1MB1ZK8Krhs7qtoq7zs
fcXwrc7LTVuc9aiZVyWewLDr/ht/4DWkVxHEQnfdhfG+iztCJngJEaDzfWhkMElWhh5GYMDeXPDa
3i72HT7r/ZQHhwR2SabV5lCc+MJOf7KV46+MaAW78RwstVJwCifLgaee5a/bx4vqxl604P+McPhh
D9gvSSd/hVA0Vmgfdo7M0mpo3DnnEcs8T6rOtQwgzj51UYX/u20tyYTANQSIJ9lklqqTN4rdELVG
k5twd0X9eXH63ubxtWez75bH6FR+71KiVkI5OGWzL0YE5kxmQ2VxchB3twxkc4+4L+dMUBxdaZ7R
e7J8KqzDCEIL3nwB2TpOnaQ2uezLRt9AGh9ySUvzRHXvjqEwGMfENiv5nvvJaKaa0EAvNEsiZ1Hj
ka+cFI5hEetmiqtU9JK++lK1FIRQ6Og5sJqWA6SpxgX4eLMx1PQTRu5zchqr8yAckAT3jv0IFcb6
6BWKtimFgUVRTSvC7Ezm2xafWjIC6QyjTLKLYhtFKjBL2fZNLe+vTMmwqfKTlwXJGV2fNzFE/GkM
HrMwjKPYyOCxdlbyJGX6ItoJ8iaz9Pe0//od9CoezfeO1GV6fLZDcQ50OEuNMWa0YLVGsl1frx7U
bStCg4BfgwxbhisNyNtljPPkwrPEcbnz/wiH57RU4NJMGUM7l5U3mX3e7tlEPhmLf1iHPgvgYtu1
7iOL4KgJVKTq1i1Wi700YpBKuhJTAnvCSKLazBQVAHCN7YHF0P7pBfdDuoCgkGYP/bd+HkywSK9U
grgOSlr/Zs530YNOmvBAUKIQOVDXQAgJs3EgtNClkHulb8Lm8XZ/N64QvydYQHn8fuzIYAVJ8RqR
16z3gqzapNy/CbPfxQvGsw2xJpx4QVs8B3hIGnQC0NXEDsUjVmyM9+K2rKq1AkXdANsd9+BSnjEn
9Dh9onkpBxtLv2RR+VlNiSxVrxm8XWXcwusODY3Xzbea+EKHm26o3b7qxXGh+gM30CzwPKI95LWT
7HQLZL+G1h66CcxVwtHZiTWxo4iB9zNuRHPJqihPD2fWDszvzNK7XJylxBikhpqZtHdTcuOOKvdt
lUIH/h/bSnTCe7Kr+dTG6VP8+Gzur/5tk94ngcuoKOpC+pi6r4dqGIWmy3l6MhFgFnEbijsKn0Sg
zUmLnyV30NoIBW98mpIhIqmfkSIwZup8I0poOZzKXdQSiB4b6uH5Jmcgdr3JjS7iQ3KbLMZl4ZMr
i3oBVpL/hSR1cV8N689dODC+OO4eGc8uaz8EnAvrvDNeTEnSoRYk8zRYtwSb0gomnlaxiwGieA3s
SjkZB8TLdMJaZP92qVIGpjSn5DVXZIJFjvQW1Ib0gj4pbWnwSg57lLrf9XQnvCzuIdon0obyMY7L
1hIOf7+cqkGAK1uctJ0xUBZ1Ks+9bhDAxFHIr4JewZ19mHf2n+fxHkv5gw/pFLxQ+ne0GCsiWSUn
l8SXmhF5PfAco/TVXFMUP5jB2WjnJLK7oo6DLLfG4+Vaht8VzBG6T4IDtrCPfSUK/avd+GFFou48
orIKyVhJsHjZBsODlNjzhOFKOid/6gGKUjhB4ED/dEW0EIWDa6kcMizw6VaoO9DsXlIrgvG9in/P
OVT7tuuMzHot451zE5aBOQhRb1fI1IezH/vIT8rQ+D7txaj4WNQkMxf96q88e/HloqNBpMoiWLst
zmdZVfvXZiuVutg2tlPGJYNRrBWiQ/zsIafj9ckm9zfGxPSgSCZuRUP1XnIlj5SQE05VHkM8VFVH
195PpW0u3JTF/jXgVSIzw5Me8nx+Bb4cx2SCpfTGUqNpYEfom1nf7h0BXIM/8B1fgRKhE97BZvWR
RtGbSZxpIvnRWuwmhb7VCouOmjqWI/l3kxUwwzwxH3imG+D0CeuiyHDbz2ILBndRQdth7O4FEqPI
P6DNGtBAaoyqY2Mv/adzPhqMYJLj1BlJPnyoJnTp5d6HDH7yKbZS80VuvtnImyPO1Ke+IpDcU9v1
yqG/Jhc6/fSlvg9rTuvjzowLoSShRkJmVF2nJHd8uXUI3wedkOj8EU7JpHsaldO7ntzcMrCq5hPF
vBvyB2AOAL7753eIVO3mXB7LrClPnEWj23kqc9Hc9s9EuA/xDTsOaw+AggNi8U7IPAWpBEWiA+At
lDCJP2WA7zG6UeG5v/UXsY+zvHHNXey+DAUdn32YDdvdbfSRSA1e9u9lRqQP5+ghF6ZLZW/GkGf/
uAmDgtDAkfASsPns43FCv3qSWeRylPgg3rxQ4Rc0b45Z7h0w6Vr6G/h612Cz3WqEvrwIfNxzMrmK
QvC0wdxc0iXycdAR0rlrv6H9+W6YetBTlrYAhb9qqtXKVO+hGquJS7PuKzaVcVTvgOoj2u0hKt9A
y+l/lH/2ZinpjwX+GbJCZ5TUACpYsEWt7SSx/Z9o/KZ3HEkQWTun52pVEEzw4LVhI1JMLLp00dnF
bxJ/uk3ha+mzZn9oIzhPy4ae80y4L2nnK+ebOlUdnr1pjrooY3j2c8XbWyZ7GH+Mw6w1sDDD/mTG
cxktm6ag22DYKKkIlEnI+M59T85H+bULOIcOE0G3ijYyCjEDapxpqBvaP4pRuaen3900CvkhsXtx
DIMhWZ8ZL7tl0X1ipYA1sdOKhYgKlwyFBMwuObI7Zcln3R0P3l2pc0CWVb/8saV9d5l2ykUm48lj
OsMc108a/4iwCQL/IHF1KBXIi5IO+yEubQH2XypUQp4FgATjaoI/7rdnUNITTmdZj02QyHcjHFow
AG6JHlacuF43RtuY+IVQQ4DDJYblO6y2u7nNfOLGyH7dyyaFb/LkfxTD2mAgwa00vz5FaOsrgIwo
PurdaGz028R5TRU9hNLSCSD4WnfF1NIJoxdAR2QXSsMsProiH65nm4xq93F+4I/G5ua2iPjNHfyC
PyPr4HFYiDZN8Vd68HHBCBCK/fa7hxLvzEMGVT+jw/6AplYngmKKvn9KCVwOf8VP80SH9TONImsi
Yj4MEYOWIcp+zkb1maylz1pQ9KqweQn+EH1Cee/VbPghjrtLZ7fnFYIX4rDsOHKOmud1Y55V55uI
RQYhwandEZVWAQeqr4R1upSjAx7KyAzCn/u6U76qzKtZ7Ko3pmbs/A+/rsj/p0vcpR2+jifGG+e8
2M9Q+ycyT/vsOKrOrrn39pu8GTUJXYD66KhQiQBGfLnj7TXgCTM9WHFZRjsYD3g0tyQqQQ2xcx0I
Ucsgu5XTJyHAyYr1PRM1CoZLVaPBciHOtD3VlBIJsltzX9vybIKvprysoE5q3BKWJBya5oFRCTlw
//gk4+HyRK3kHG3F0K0rhA8uijDUpPM5J3LO9VXkvYqEBot5YsdVJ6rK+EOCMzKgKwq0idl7pSGS
R3cWKnaZLfCWAJ6DMyTtBA0Qee8skLnUEoQt78VmOTpsGZ6CeyeujR43HWXlwRFtIYYq5U4pm2FK
Ez1TMBSh7hYacjA3j8b0/VrjnYACchZ3HakyZMNdz4PQZhuxCXeZiSkF2P06FAxgAGfCRq7M9J2X
41r9Y8S8DTfoJkSKOsOtob4YdEYiJz0TLgq2uRD1uMxc3wYVgpwOOyhmLdq9H4SZOGRsIbjzVQ/S
+1+m9E8ng14JgBcZtj23e2kMJ/nFkrHq5vRUxC8/6kkq1VaS/xEhDsvrh33zy83NmCXH3R0c/Pu6
FVhIDYIKAAymKVzx3BONssjNH2NiI4/8NH5qjktFiFIH9/zJjqgAdkGdPQHTNqlMWd6nmB/4Ddv4
V0vb9YsgEhr4Hz38PYQrKJd/Fi+4oDl2uwWVw3zpKtwMMSzZBbZ9f9W+JoqJISs1NZSKhzjyi3/+
JPzr0CzxdEX65nzpXebatl6iBfMxmwF2D6fTQ96FNvRA2aEQQ89rbI+jwCRJuckCpVGIbbyJ5g50
c1bMWVXxh15qsJfwEbkEKV++rN3eEkpC8NY/9ibwai+hiI9VooetUHSlSQH0ztDls3Iy4fCiO8Gd
b0iePnAblQpZaYBFFApQbqv/rWd+VxCe7M1i+ntcJwRzYE5RwscvMK06qVNMdvSdK8AF9ALTfXXt
PwDIstX1fYYuvHn5cc2fW1THgUbo1BAF6B/wmW+gaLviZGNBdxeT+jm+asdp/3s38fwtvUj8ZUo/
5Co2+BSB/0RveY5o1A0shjrs6jpM3X13qWDjJtmeABm855S6SkJdy+RFDc+fPnspHH2JIPXchwDb
UuS8QCpkNAvmB4q0MhgcTlr1kAcHF6Oudf6qwpXOK4mcQO6Aa2tdANmSm9eaNqkEOriKqWeynhU1
vFDnEnEDM3evNs2x5oRq1dk/fBGw9RGuKjMoTj8uS/0/q4Hz2YOrmOX2qp1ZhHiJ5xeL7272K/3D
p6GwvWB4uarsyBU04sy8ikKtW/Qwhjl8BhwZxoXCUmnRAmNguuh2SJIVUcZx6qSm5cW/xXm1/TZ1
3bEGLq3lAuCwLurAIUgCx1QKvwCw0kllWFr68lxvIX/cdud9cdjzKk9fBpxTk7YhZWGabq2nYIEO
IK1e1j96PYkNCCucW0Idv2VS0gy4vDsgvG1p/aHCtLHoQb1QXHjYBdzhSN+vtYcrdqNGCmImucOa
BQsEA/MtZ+U62koDx219JDnmR35y44jj2hPNrSdJCHJS9IDhFfA3XiD43GWL6CLoPndnkzjxT9YG
xbpxwI+G/dJW9few6oTm6M4qtvZR2D/e2UBR3ObwJYGWHOzj9X+O5u3kRORUG68nXyVuaVxUpPmZ
fY1APdX810Yb0YvMckXifbvn7PSGfdBwtBPbjgKUnA23FVjNxjS9ceXmtt3PDXNvlCgmIrZM4Ewh
Z7rNmT5SEj3aVr660owfJPgmz94ecOdQ3O61eP9kKxHHfEcCAKpoj8y+UdEbXQSdToxeoa9myaUr
aQEr+CUaAl71qL8hdp7jQTD0xEOfkFFd+c/KJIkaY+fbC5OKO/83klUGZCPPVmYvyK+s09wawTVK
M46w4l9MxaKVxaWhN0njip6UHzThEWG8P8+JSu+8Brgtuayc+8skcqAxKI7UtDOvNHbHpOpf6lAW
OKD05KxalefwL2h6gWkMC11qepVIZVHSJnTwPoEPJJsFbOw+6KetOc4Ayte4F6EJO87R6zk3rxE3
zTzZg0Edq+FlTLuNBsKY7zkZSpJNtg3E3EAZpGmJ6V+ZqNI5R1eZH6cu4qcfXe91RPvbEQKZ9gvL
9o2BxtimURGnmzpuT6yM2oSViRmxB8tI7QaRwbBQNuwnqheitg4Ifz27VvYcTSd1x0GrOfWe9xyp
cuxA5ug4X3k5v4RTq7d6vgaB8SM3gmk1h8TuAQtglWEVCTPw7OOb3uap0ZJXKLcvujW0MtHxbHYi
FuG/884JEE9etrSR4/Hhs7Pxa4LOcpZhIV56xRoLFG1uQex85TaOHXFuO+6vXCMP7beCioBIjwWV
eUVeEf3CUSNEZfN6Sa0fCHTRvU38HNjHezfoPvvG7C01lLBfLqcxonhMBgPlrOdozWcGE8cww30n
5rXiKuiXdN+LZSuqASfcvMU2Ck5qGlSISG81b8HhEm4fybInUBkBPhwp8OJkN4gM5hCbjSjSbwID
rAhR4z4XHv2VljiSM77Wn8XCdYNgXbEsjurbSqhzZZpW39lBf+SHurAJtNAYWdlMDfBXcCLOw/pg
vQWvqS7EvtQrPNyiw56cFEUkMiitvM/hpgXiCQDohM3boZ7LH//WwlQm1GvrucTnu8atqGxBoyw5
sFQx/d2koGVXbgxLAAmiDKmW60x5IcETN8kOPxtQUeN7nwHhgJtWBZKuY9I5SiE3kTofOC+rAqcK
a96uHGn+T9i0TJwnFE5HVtwdPkR3tu1EfNDrsrnXNUQq3RV7nrAdaeZrphvv7zvBLbkjbHaPZ4w8
uhT9ZCWc9vP1bhBWmtSmmW8UQBxPWyBsSQq5ywPfuHbf8uOff98kZWwJgLBQTGNk2pHfStvuBYwW
v+bl7jLl+JaKFscjSw9GxW7IcMJa+g45kXGD9kVOs3Mpotd/CBUXAFUs+WHwvui2WjiJvU8l2M9M
1T0AbkusLrWK0//XzRd86lRoh0RM0d9Tfoz+dOnCLo7oI/EPnilTfRgtolpV/Xf//lmn3yM//zWT
2t3JO628in0Uxj3h9wFtwPnxL5LZ8T7PsRU9a4dwdNFrI8BiP8QHYS0MTrLzVKvLZk/WWllvAUkW
6VzU0vbpwmrq56/gFMVn8kSiCtJ5GGgsIzh52xMyF4UScls5iPNAD4UPK6RWbdKEQo7Sa0Kg/Bje
L4vSrxttw8vFF9C1dGMfN8d/O2lwdnrp4X0TlT36ELEO6zpW41o8iw6ojTiTyNE54QtWij9Nmim/
WsYWVCSiClxn8aTSH0Xv4wl14W6q03YcQdzufLhyrGeSHv5J0F21+RVmMLm/ImDBg0l/+KubRYSq
XJmCBZ26j6XZWu4Now77tewsuWL5ySMctw2YL0VmEfgQN96uoVSm0sm9sc2EdZCuE6YNf3XFHS2S
1vkhO68bqWC0JnY9GNdpY/GdnWxQ6Yw/U7mfomlhEap9MckvSbzHeuyxgxTF7AUk412M2ItyMlMl
DI/fk2O9Bfc/ql9wVtZhYqSPCp12ucYtkTxv9tfVnbt3Y/gdprLVLfWu9D1hvd4wX88RJkGhaJrF
+5sYHzlvGDzSqRxqkpoNrlJlEPvaeyavFpJauQh6llRg5AQWslIUst8ei86dKXRaciWVT3z3J2wx
KBv7gq+nDdyyI0gTLFp45LsHXo0kZtl4J4782eXcIYkSrOSiGoz7d6exbcTeVY9FgzENwx8JMv1n
TeQe8eIUGnDDuc+vr8ayGx0L8jMXqpKc534iC0FtrTkpAzKEgzyO7TNAfOTF4NXgitikehoKahrr
kpPjMU8PYHFIVgJr0Im53cxsZZ0K/8UgYE73xFnWhz+322O57EfWdg9LeR46qVqjbHMgK2fW1aNg
DuoW7B0y3nF7aOtXRSXXC6kzWUDY2KCSyOsY68AzkQiKkmgERpMm+5XfkYkluYw2dVpuRh+w3THk
oL+59AYoaBQTHWuI0yiIUg/hcSc1nvGzaf62Lyda7eYt8UvpRFSya6gKf9VaGLuj4enIh5ytuFZV
TnkRcQOZN5xYeCYOm49wIJ8fLWqZqTR2kAe5A/llxb+he1G7ZdeqwIg2xNUfnL1bSncgmoZ6V+oQ
nuCtmKhRRG0ARB+FcKuUDB9484i4G1zH7ZFegw5pWC45ACl+T7/E3RWmfTtcW9ltgamnhsYOhzbK
dROooE/f7M+O5OKJ4z8d8E3qJOdqn73HP6oyRj8dG3A7CkZz82VUxS2+pdkcPEyGbool84sSo5Pg
mwq5K55JtaN8+TH/xWM86/rAzrtLpVFL5mMzZmA2pdYXxLr7XUzHFUw6cJBRLKF6iZAJNjh3qqNa
WBqx6StD0msJFZwCMpYYdgmQukv/X3n8s1FGT2b0wEIq7J1rwudXUkqgmX/23NNMu29PJioUzQH+
MUsp4Q2Oo2IHgeCetrvt4YnvQmA8YoVCCuCFr8sM0qsQF9LK/9UtqmGv01KDDVqrvKUHU+3ee1Gw
bLl/VqP09Drjlquqd++4qPIAjcxxT6loc74QUFR23v/Ygt6fqQ+qHCdH4Bbc3S8DwQIuoCtrTrUT
ChNlbSUve5y69VPERN/Yxg8yK4PUsheByMyIqZui1ljGcjlpHWgCzK2+GgX6cmht5EeA2nXdVZAy
YjdoOfX9XTJlRM5kC38nibDdpChHl7MekUB1+2pnNBiKSftGOqVk6PIJoOsmNndRpauYgJvhppUu
32RujeDzidcjRQDKyMc0OiusjpPSrHMb1hiBZUYIR0WFWeughpgqg6ZDxoRNM8cHYwTHJYPLGjfb
r4v5HdjPAIW0R52MDWusTB68S1SQQ5TYyYKUwQ9sTqFwDEcNhITQkHeuV5kcsOwVUXHwG8TIKelO
8Dmd5sRqC34Yn/pSdzv0gQ8qBjojGTqYZEUSzmK2MvxbhCVW/bYEaqDNqqWJkdK6KcZ+Y/5E+hAa
QTZRf/U+uR1O90g+4zyyl8KGeC6VfqhpP6fdsvBPKd6aDNteFL2jubItFKvwFnyl/hkkw3wm2gKM
ACvANhjYKUPeLqgpNpCXfD5wkfmS2wgxU0GJ41xyFmeLLeHns3UQxbGEtLd8rJYsBKhNRH266XpH
y180iWNq2Td4eeaHDF3XBjAn59rcnTU9Y7WE02TZ8K5atAbIe4/U3uZlMdqziibkx9RhRDoScaYw
/sLUS1G+m7xU6BtR1j95es8GSNgJ4nVH3IAHn36+rcoobEPX3EShxWsUiXlOVO7t0/IsILXZYy4B
zUYVN4ImCzdZEQRbxeHBqUE20sILX9nTNR6gU7m4MVv91SU0jCUKI0F8LTuujgFZSsubidoKeGxq
CW0ByTp1SQ7hm6L+sRZfeTyFM/P+YXtucWhJUdxhLHjm244oboRFoUf/X3ObWKvDocYqJtTR9KE+
ks0sB+bB843UjwObgaLQiKkqngAvYYdfKxrfOq2v82MvVX25sk02Sv6697qBJI4jvMAuhmjGi9aR
U1I1jkNOyBNubmCXT0Vr6KbYRQ2uD3AHhWmS/SFw2LzSpazFpiBB3qDFrlFpBI6PcVVReCRsRhf1
aYorrnolaG7uBLZRrmJg6Q9EjhlABG+qdiDR90lC4JblzMbwoXi9cgBzM59J0Hm4sjCQqTxBaniv
JD54RDS03a7LrTbFSqTyVvtj7HArggPA+i9Ft2ghhEbBO+FiYQ8sTOqJdBscZPsAZpz8zyJdrUQJ
9hSI1ymL0RJj+IBqrWzoWLw7aOyXc/SZVwboySCHQWM0QMOYmqvD+fCVf8nacEORP1Zbg138fziL
ZpMOr3Xrt3XiQBjrsJ2RMxu9x9qyvJoz87iFrtI1h5fxUG2ArOIjqhxz6ESTpXaQXSXReTVgUins
YrX1mDjabr6jBhACpdFk/15rT95sE+rbvahquEH3wfjOU0bJMGci+pHo5axU33QI3y5P0DEstuyK
AxO2wUbsVBz3t8n1Yyb3VL9p1EJI7YdSD9xSzDQqjz7niYP0fj9Q7/KG9R93NdQyi3YIjDjwCjNY
t7g/Q5hTcylUk6iVbB9+awLDiFWrTAWqkyxvhAUiOJeNoRpyepZZHXzr7IpwqexYxbOpDHJAXE0U
bIgMHrN3i+2hCi7ZTiuBStw2LMV3rVbO/suvrERN8mz49x68Nb4au9qM1BnossSPI7tdEq1reSSG
7/e6hrzNemF7yI+vRFvdghD8HZf+GSEqqwarRijorCm5J/n8MoqknP4zbAfIZKJghkNKl2P9qoKV
Cn96I7eUhiR8Qm7AGx/+wNvRyloKtTW7t6whQ6RMTMtUzo5xK6ub0VQ2/SVJgrrD7frXMVTpQlZ/
L6Nx4VH86Y3Aty0ORIdl4n+XniDmLMVLFSGF0K2Qcjxl7GWklTntjQAs/yYSx5kb+mPBOrHQGzL/
15xKhycpzY0/q8fCoddcJMi5zntWFKUilC69TwQwfxzUbo9M5pP7yE5qBx65116yT+E509r5xB0u
+BCHBKDLrRb7zAtz5wj0nbutpaLXVgInyUXAL38hiLJqig7H9eQl3X73wYw8PusEEvhR05qkLC+g
bgUAVKj02w8IKAWDyntHka8/fJq/v4ZfW9BtEaqeBkEd96LMcAbpw50qOsgKTNiJacuEBJoxuZhj
nQ9/wrauA6hZ2bNw8A8VD8sFFM7o9RcvX8V3fDZ4FhezEpuLrj0zvmn5sEU8hBabQF3XXK0q5oZ6
g+0WWFstEpIdQB6KqcfvZiePbTb1pSDlTZNlCq6MnCpxleQ447j1j8M6wSb0dxBmYN9BIDrG4T4u
/K9XqJ4RqqCe+Bm7qxbD+YVADLeRAZU8ULOK3YvMOzMRE9Ji6S1Ls0Qg48nOWHA5oEcHkuLguwPY
FG748ENkJWz8A8J4TUUXxeTUJlV8HqyvR0JIwQ+eMD/nasXR+UVPhUzZgq2XEVDo1JPwSRKUZD/D
Y3AEUCuAQx0UwCjjH4pDLIfMHF0ripNFhLlHrMFur8I5ojDBxsczpxU57ZWq7LrFbSsyHsUQUvNU
IUhm3B7l465mBoYlR/B4SLPG3NLLoLh+X+Cso9cpI53Jv1i8aJf5cawDad1rS9dJ6cdsXmUnqngt
ErdluQoYRDJ6ZmsfZklhEJS4mTSFDruUYgAFn1Xpv5wpQx1+IBOGqswJXmTL5KP1xS6taOj9sjrK
zbzavaODZbd7AQViWLkg8BdGR0StaMK8Q6suv4Q3hulqwN/j3Pd71QQdz42wk+a3+ILqnrgDmuNu
rlLWcRkYKCoRabDDzPLcvimIeGHmmHUhb/JpIhSxSEqikK6VRV3lG7lg+ZS0xk67Fby1UFfeOs4m
rpQxZR5dBA7oGxd0MAnWoOAHs9U90DiWVemHQIrZFTzFBNCA2KcBz6hrPyutAXG+cUr2AnfC9PNQ
/ZZibhXVLYal+uBMHaaVg0MUZ6KtQfJXyDL7JNeZZR0NfsbXF5Pym9EYvR48czdSKeaWa6oqb2xd
lZBwo1fWRf3l+Ri9WZMVdeKN51chh5ivzmKNxsSfmOng4c2RdzCfFzULM7BjsCyg3z0SH6ktvVNC
QzweO4GscK/IVUdMFQYyzh86CnpDzgGTVBph91dXFOC0syRhdc9oGPwckHIJI3R9uTvax5AHPizY
zuAaGECC/2vRlisyY0oHyQNCq3Cy/l6ZtlDZvyrSne6jopVWzrYuIJ/j9gg3mzrlgo2BSvugIQtu
z/uiqrf4KLwgHKMFePa5dIzCyaWmzSbN2YcQy9/sVOANiCQlGIptLKrfxFlgQaS6j5m9Bonlsxg0
B+ukJYyIdo/vfrOzhR4BHjuRHSBjuKTjTgFo86/yFbSuuVukWtqWr+y3nzAMaabVjgp0/1azBJs8
cJ5e8KXVpgdZ9kkPfixop5kIUP/rEzmRMpdUnOBsfzH4RchPEBtSm8Iu/9C+Xdd56v+L7v2UjFHj
JtIVrhCJoRDAgtOe2Q0PMFrEGJmeNiBuvRQ2Jlu2EQmT+cDppbc1gn/LrYk6/Pg5z4K5/Et12KvO
L6rei9jpHWft7SoHlt19Ms5qlot6LIPiXMRKvdzidgqIrYlBAfUVMV2bWvePISjejRkCV6OxCmKJ
r8EkgGABY2Jm+xyAGJKnhduHZ1tiqCibTHSCDFhEk18tV3ypVrH70H/ZfbnTItZ+fDNZzDbyyLFV
owmGZJvR8eUI86kd7fZYfCMaTUPz3CHN+YcruLqU/3VOpz9aarnEqjW4Q1cF+UTrdqTg6R4JSMsu
PxilgZ2aaphrpag55m0cBSJyO0fv6QGGbXxYc26KkXeJCEZsYDbKlpcRQDeTy5vBiKd7tehFTAfc
hEu3KNzwOKExofIQQvzgVeVgHk4l6YJOv4reqWu2khhuE3+NRFvre4W+9QMAnX2lnBWuzfbPWfsp
5Yh3bkPwMBaRf3ZJ7uQ5JAYIh3kpIAd4uKXJAItv8BJJELXrlAlKYJjskJvOIpAq6Y+0qeHGts1E
T/PxZikdHaErje7VoDZWXIuY53vDtxp10T1u8qcZb1MVEvD7heZmkhoZuKbFRZj8PIe1sRUz+QCi
r5W8GfQ4KBLdCU84A6Rm/GNUpJSmCNXfrLyKtYaWas6A2KZOmMEoeZCNr8l11qgG4L4WAS8veDmn
EE7hR5xotF07r1z8Wt6XFc1ZhUMqwJfqlsBizUa/UiERP9BNrJhXXY5pkPw1noW34OUjSN0r6drN
lBM2tuj7f0LWb9C+pFcoBO5fkN1OlLox4GHr6g8mt78ZlUbb7oI0KiASFas3qKdxgBSGGf9IiyEe
/kSIbi3Vz+49lXqCbHq9zymZzjD7Sjsuul32rx7EgBAHcPsoGdmMTPJJkEfmgBbJryPP89IMHUXb
GxM1Rw5sYjZfakF9a9wWjNzwx18qnOeEHiolJi76tMrgHL0MSeCOK6tnmIedW4W0VvZx/+OMsToV
X88UDL3ky0HuZtyUcVYB6BHFIIu+oaV0wzT0iZslHjF8rJh0/+seVqJxFkNaxKhmL7Ev8RHpEai9
9z25tRxdjmuVF+/M82Olbr4YT0gqY58uiuqapGW52dCWpQKKQI6KGvXu3MAV89ZY03mdYmK+XPbl
BFxVG3jL64bCaAK1sJArDYNV1lJwhsVruJ13qbjyRP5s73goA9KliEXEFndf7cb/PhACVL4tcIQB
b59PvX7Ml4c+MOM0CczhhBMVq/2zkDJhPMG7+njbw6/dfPR4v0bC+6IhMMykiqtDO3MOOCz5vkC+
+22a6JP3h35CKFIh6Ps/EnlVlziGVMlZISy54+64Vi1sqVnxcNytTsRc1c7UM5wDu7ldEm0oX8/S
JSZVhoHFLDY7os1JH/V5SJV7/EV1pt6Jo5nF8wMfLLF/7m7TXPwOUt1rVOH3zf6IuVj6v9jxFxKt
2rdu7x5tlhLPSZp6oOtL/K1URB1nkfskfTfcKczetiKGLck06rAQhND2Env3snDNKewJBnPUYSVg
imjKdBQxIbfipnhYVECOGAK7VXdMjWWM+S/oFHR9KZ2GckWD7c267m0UR2swD6ohdC8uCh6PBPGp
vNzmhacRkCS6g11Pp3PBEODQrWaxsAwRyZp78BZfG/6TGLZk+slKVH8MDQXo1OwluRjpvE0DPC+l
KX55As5skrHmV6kwNkhcnlt1eSPXnLjQMsYhfLS+0O7RTOIBPMhhhH8jeWCPnqXQgLq3AkMwYzwR
5iA7QU7PfqZRLPI2IBnBXo+ok7nqogPOoljxzcOd4M/kQC1gxlbyxyRKYiykeqLy7LdKW5FdHsOb
7Xz6+D98ukr5OmMvJ2PYpYByDQxU6/mRBmsmJA3cWn4oYKvtDu2j1jW6lCpiVxQwPKNXnW6/ewMx
RroRNS42MN0DyxijQ74mRAv1oy5vcf2ciEq0W8ostrICDFkkMEJr/Ov3lypg4MGTsZZHEv5sCDi0
KVKQMUuEpaJFleLPew5UJOi4Agj0W2JwMcO6gaHsAemiz1wOiskkha3kWAJHCi8qCdxf+sLSTZns
0c00CDA4hpOAWZKFwKcAXgJyUS68IlqaR9djYccTFLgwerT1bG7EWwPNBKa397D6EGgOWoXBO9pG
NbNTE1jaXPQi4scNyURlZzx+fX2npUxRnIasU9Wy3aQncE3n1LmRI6/CRlrZzkTVxY2LYq69nePZ
87OwhiOtl43k6hVMZHloylSLF2rhGbVsyIkKg+ip3WsVG1YM68sBjJUY/436skckvEOltiwTtE2S
XRdOTVUnel51D1uRbj4AtE/XtokNgLwuHb0HBwf6TBSdR5o/wJ0cdBBTKF8v6Vw7Oj3M8+HQSzW6
ph+EYSR91cbMOKhbQ3Ci09mj/s3hzPnRKGYCxIckcZt6gHpQ5m9+EURMwtFlRWsCNj6CzgS8omjh
2qbQXjmYhTU63pdVfKQ1GlHm1Xnf+Hd9OAlDz9cLPJ5l+6Wxgl/b2kSkIEI8SmKTDaa3i86DFp92
ui2K1DOChNI4n81LNVB2Lw9xgYosHvrJznSHY5TbYuA85W3A49HeGH2h4nPfK+6rZh+QfV1xXc7m
z0PYqE6ePnMaeSYHs/S4uWwzGZkia3/DrOTEwRGIJPSBKO40nXM0jsgyVKmKjlvlY+8qjQkfw2dy
ydwIrFTsoz4ULtBh0pE9Py5PX2CHhACjK2TzpXOllDtjfC9OCHOwHKekeAvue7FfbOve+MiTErvy
DlNeb1yoPSpao8RQZ2xcRmEBItgDhsqSTld+1F54NA7ZxSt81K2wdunaAfoBKzRzwpIbyU3mQB65
VCKzid11PyyhYSavikTNQZSM14fM3qgAXAlM4y5QcXkln+HGZoHicLMxSPrviYpC2JK7ppvKF/jo
SHZEwhkFn/tVNeKfYBdJPO1IThTU7l60TXUJ/TnnjrGm3eSZ46PEqIjHUfL4xNG1XOtno+XtjimJ
bpof44ZScdpJewRmnUpcjA+TYg7UK0OA3sofxB7PpnDRrE34GCOaFyRfFnJOGvnKxGUjhW0w6UFe
sRLP3W7jpVo+BZcPQxcMhQbFpGqi5BiGqqNW/6MSAixcWSBQY3DA4R9h2c+mDRotpVBao2onzyS3
9zM40zmynGmvRd5A/x3QDNuX8riNNMCpQbCb/2jT2Napb8WWoj6EnKFID0DwjgWdIucRg9KzzmWQ
e1utbVVuyLLYlooOc5zAAIeOkUj8ITmeKEGG5pbUN69s+P0XU8eWoOOuQkqneZWgBcS5yB5S3uM9
Tt3B3LmOmIqDNRGUYnlaMa7mmX3QBpmucEWlP8GEa52KXgY7Q8gDkzi9a5ehQk107Nnf2s91Ac8v
0mNK28jGAxqWN53N/go4ehur51PYfIc8XAyYurKlSYnKhImFWStGL1vMCBNvtOkjk3cKe50nl/14
dbn7LDg3RVV4e/aO8RAR49Zs27y8wQ5Wb22Cr7M0kk1CiVfU4TiMVSPEhEFOKa1Zi1jwtOMXbPYf
9ywTtRAEyNmES93gN6P98GvI0wMlapbifyXLYS7E3//oCeMx3DfUiVx5KArFd/O9l/JW4vnyLHVd
RDO0VuL0O2cnl+QG4cdQ2IloSexoYbO6clUupmD2uY7XU9vpJy69MLBGU2Gpye3uRb9gfGcqKkGO
mBdehE8Li4I1lIK+LymbfboODHskagpe5F2h63/AZkc4anuM/R3ZHI6iWedEPhk9UI3KM+OXuK2A
Gs5sILFiBSl3fq1F8iISv4i4sd4VPugtE++1adVdJo26Wnwr4lTQLc4JYz/8QOitUlczVPVivTms
UMVwAmlljpl0JO9J49WG2OgmSHeNWC9yGiFOxkxPy1L6Qc1XPQA/EMr1uMTVMfMgBCMz3jYL1bIG
zsPuL0WjYyVje5dVXI/SwEY1Cky6dlmd9nFAVd4Pbhfn74EuMX69rrMY6DO/ewK+rVKYic9+AfHp
qOrdj6rVgpfOuJHPxJe87HJvXG3PloKSOcLb3xwxcdUFWrCJWnb3LRpEDvlwBCczHe7YYcuF4Lg3
Zf65hDs676BdJRrG0gm68OM2hhC2fdq0ZBX+gr8/6DmD8ZMRuXtNzeftvH2kxvpxmsZjChCOpfAQ
4Dq7vwwmmWf6xrkSjcFQ41pR9G2gSEZmnK/CPgzagrs7yXkwff9Fkxh8wugIUapbE3xeELhDWFQU
A2mNhVFDZpMVDYHsrYIcoWtg7N8Og7RaASVXqWmGuEi1g9bHRiIWeBoX1WtBcZ2JbNPxqiaHeRuh
mg3LgAyUWQo3uW0UAD8P4S76DWRrbphhPpOTAB38SK41NEfdp2wWdKUOtSfD8HnGfDe4+AK5OjaS
Kjs5WhEnDzTytxR7oijFQ+y7Uq1mLQr8jwBcAxKWoFPVtJq0tHMG49Bqo6zBd+XwgZ7t0CqskVTj
x9enfsd+ffwO3HpfQjSrozoDkndokJWcxCkIH8E4+RVU6VUJPKaE0MhOYeU80yJEAU9Pfm13nRPJ
/Y58zH7JUQZQmFXZe6ePzRuP58yBdP+vxpt8w2qMXV5YGp1d0FcRQhSD0moFdHvEtYLMomqCFKQe
sCvWMco1Ge5/Dw9uKCu/ww1aOHUTpsMjGq7g2E7MRzxhS6Ni9jx6t/8s1OMHgnxr3ysJUdj+p0x5
fbgVvks5tL9r418P38HSUlSyNk4qbcffF0i/KshaUrciq+Fsah7Hb52t0zMF3QnDvJkyJ6tVHwRR
SBwuGD60fVWZZrJMnXdGres092sS2snfB4u6p32pAA3zhiKl7vkerVYMlXIWmQLsVrom+fkdVXC6
VOg+HiWwpaQGGk1SKMn+5nnENleuCUDCBlaUIjAxDJpmoWV+b312fPL78wBclyyskIcZoRWvy2d2
5GJmyntQ8sfqtvKOLB45M8W+ruBqXX7ryxzwIuxWroEUzjkCamfb9bNXIWCXAqoV0gWVeRMlhHQl
DQemnSZcRXhrgZ0pSQiH6nDR/uDmUWIWMUm85yzUjUd9HzREDeGmdOmAbolROQQ+/Usf7DfnWdLK
czlgtCbeUvDgkWtlnazs5Kyr7qhu3jgviV7iHfXWv4JxwQJR0u82w92dacqn58g114MWumi055i0
3a6pTstIxiVlazc5jZRv5VVDYQx/xr6C9RDQkqmRmuy5KT4l3aO7Dyxvpf07t+OFhYFbL9sscMmD
wIJdHtAJWGkCRavh5GWjdhjl/thk68TyybpltpuFqWYT76/IEknyVG96mUCc+9wqdAfaHlELCXo3
AKZIDxs8AfnotF0oNwD+8+GfJCigKMyAjPTRuxm581LPYsYxhBlQp28YIVx23Rgz69N+rUhhDeg1
51wfr2tjfSBA1HKq6d7wIVcpO8gf+a8CcZA2hmg38hw5S5jOoAN1o875PQteo3+kdzmEipwwgOAP
sdNtHYL9JwGVcRqsVITt4aL+9/KKr+7OV1/9ipqTGJ1uwyckFGf+vetjc+eUzuNDHi7t4Wscvf1Y
4aC9PeJyVccwICaOvB4KDg2lQn8gOCXEGpCbTw4XPQJdmg30QMzz4yBSEAe7ECA0cdJRdjLebJz/
3fHYn86ZGx3+yNWiWJWjR/ky8yo27PnbbV3b9ZC797dc0jGkw8cpP4W3hVLM2a97vQcxeLmvVBnu
SpefgkrKS3tP8kbIMR81eJZTYUHTb6sCRoDJQZEq5ZWrTiukblaSNpasaTHWUmL3IVv0RBJNIygr
X3ZNXDQ5FP73RKaRf13mGeYhF3MW4PSvsp1+SjCieItDddICZNYTzD/vC0mLjaVk5GM4cbUeDJeJ
9kFvMKVzwr4EEYuLVnQcVEaNw2NxASYj22RmuQ1vnXColA8WOPk6CTb6gqW6wJ8m0GN0o0G/+rcU
oAWu7G8U1wGjjhVxW3I+kg8w89jt14eMC1eDq2WVXtz8lkdV4CmFiA9gPZEhxHJxNebYLM1YIWJe
qJ2WKMpPcldjzCWmVRRMUnR2XquC8ytOkEjPuBuA0XSMf85NXMqkA8xB1Yqiozuz+7+9iGjwPXgP
DN9Eltya/bmJ4TvKcKCuYVOYR/+8ZTZQgap0wDbwC5YRwRPwktNk+qfpGKzfM4QJJqfi+xCijID7
hYn2zbXVQ03Ibd0OPa4V1MfZH5+Si0UAfWRjIfVqpvH0gixFG8ID2Ysool7shnuweSSp20Q9+c62
Y2R7dm5FT8XQ+c0HdELEZ3V7vejpiLZB37vNi6DHAUhoXPWUatfcwrDwKwLnqn/5GiRZ/sj5NHJB
X3EzOXKeqLKGAYuxmN2BxvqE/EZ1+azESXyiSWVR1CX9vsz55AuyB2eBvUyNNxS1XfDeSQFSElLu
INWBeYYA961ecmszhQcvdjKj8OEO2wZUHq0SZY57ondU/aNdBI3RxTVwAIodF8C4P8bGg+5gQaBo
zSo2z2/cY+eMCBEb+lw7rDgf4jqR72mCdmTTZPEUvxEn7qbBNRenuITGJ1vNDWIgjM43KagDsolj
sgFFCafLExKzqDtvunspQE4vDxPswCCM1jjguiyDX+mTFxnQH308Bcna2c3hlLixEel44vO01rGb
mZgHUgs9x81CB9AH8tqMCx8X9t9UcGuTlb2NASUvDWgIQZ491WDDQGJVAi2ztekseerWFSlL6EJq
XNNn/Dncr7Y/apDOW1XCef15J0aAHeBJEUlaF1S8aGZY+1qRl1m0W5kD8r5qxmklgNOEA+LnelUA
UDlDuPbJdvG0V8u8EXxKetwIGVveLrJ+I1Az1d/7KzdJA0jQxEJ9Y7Ui6QXf8wuayKRvRvggkm9h
XOJOmDb/7Z5CYXBPuXpUj0a6w1t811n3XLIO2RnxA0Lhh9JyUzbrslQU9Ie8xV7M9JFwbRK/Z9u6
p1EbkIsrlCdoR24RFnqzZzVuBUv+FwDSv/uy/H08TqoVQntwsjZxu9ylFUh84FN0NPEMAR6qk6IX
Xm8Zqq1IsbX13dqBp1eIlkL3TRC+J8elzLuRjBa4YPwgD0Q8ohal7znjYewnh5tlwgkx7f5lalIs
RCk+bJsXd3dRC2VTEc2Swt4jQjsQK8TsE0pOiOeJOvXXNEzyvDq3GEWwq1R/VNIBB/1kwuOKvaXH
ApvhFgIWxz3/qQ6CTiEBtaeLzMi36pmT/gY21Ulxl7P9E5qVDchxdIg4Yye/Vhbwrhm2ISVWHt3s
XkQjqHYh6WK3ggwyyTjDY29smaFHTiYTV0FcXX3WusTWkiLo6SpHjGIzJbguEjGqBVB7xysZkqhz
hYdkPsYXN55asQsqrZumDx04/y5hcGRswdBBFbPkbCQXMdwwCFXUwds/I2caM6yJVlV6LDX6bC1m
MolU7dMbPzgj19Teu+Ksg1en721e/1rlMyqBTdHky8F81Dyi5699c6NQD3mbHgvKtCqTeUG9VjH4
x1NeIIbB3BQovWKx7qK0oS2BpAkAH8jbSGYg6MEDBFbsQP1Ec0osRXwEBaXUoGidehz7kVkXtutd
MZLqR+2JwLe3Z3nHcUVxkIj7va7gypelvYM2ZzFg2Q38TU6rWi66eb2QVVyxiY5PmaB0ptjXR58Y
SBcCpVa3NgQYdc0pEXWrTHt2Gv96zoX/J7TYf7d5uy+ZMS9J+G9EcimIqSW9mTlFKIN7/CWsLpkx
6BXiRVYSpmgWfAHxp4FVZRzSovkv6Vh4mqEnj7H1JMqFLk1hQJrb8+XtvnghE0dvDhJFAuLjyTTr
JCI7rbNvYp8r10so9r4dd8GiVBQKNvIsjMNcZqFN0TLgw+hfgXs3OALk8cC8bsT0tZfbZsr+NZsa
z1niNAloVM64zs7SDGc/Ayj1nJwiEwX8M+g/iUrWRi2/thv2rBeZwI48fasBtlNsaoTihfNoOfjh
OszIdcnQAJFoaLa4hYd/qhbgDChEBKLlaf1tH1/KmPGBw5BNCSjqdnKsb6KUVC14mW4vT7dgSb9K
rjJEpkPSDLHN/uOVOD78pu8YKy15VnTudgN7ANN4I3kTkhp4uGfy5p0G9z6GQxyZ+8NeJLVcV3Vt
Up1Zqg/3DzPL0Gr3NooNdXxIqXzN+Ux08EgbRPDbEqJOsWBQ5o7UajM9snni7/iiolfv3l9LgqJp
tq3s5xDCxfriuoU+kfPnh3jLea51h/ijyDN9XJ0ozzMRNwcGREvGvYZvrQc/fL3AXmav9rkiCVFF
oWRnxJbl4jp2UGYh7WgWjrDfap/noRzWOeCxx+jUi06+FlUA5HG15PVGc8vR0fD4tk+joEjgbBip
WHj8QG2rp4/NJ6Cs/f09ukqUT7ZVGk6+vH4+5C6Xu4FiVh8FoUxtEJRXOWvM6ZBz7wZ4S7ig9bsq
eJGrxrswb4tzGequFXiNPMfQp4but6bha8ExnQ6pD1sSUH8JDVKFiediL/efpXw6OgGGnLvjpyHq
bXISsTNBU4fo//VYvDmrZsgdfUN0RK2NB4iL8AoNOscTOIZD4xOH9CibYJUZdlPe+/Okt179ZwWK
5T1ynycUzlbnv3A9iIRVjhHTHndoVi70w2ArKd0r0TOaOQE6nKFRCc1lkfdWTgoylWss3dy6dcnQ
b7YpjMC0WVK4+OL21wxPNWmE4Jg0KQSevMVUaxm39XJ3/o15AoAy7jKIX4Wq2/h0BRrgkdYHaqnQ
PY5F7aOQoRZJr8khyxdhlZOLnRZqB2rPiMkYsHngz+BDpplAK2ITzlCEBWuaF3rrAHj8ms5FgaIE
H6FdWJV8laP2BYsA+WQCTBSjgfLKd6TVGItOM2F+ArudAvFHVeOABs46wu6jojf2wOMdppGiS/u2
eaPmCZO0QzooyEWUJrsqVRZWGgI2CsdUcheFkXJJ7DuNo4nUJEzq01B8xeT7qQLy5rqCzTgbGXeY
sSu566zlrcMbnZcJple9Kv282bQjuRCQIf7d41dTo/tu4IPLviyDiWnCSFQLtw2kdXM4EMWY4Gl8
qCoauXFK8GLjMzgxYbTsJ6DeoqNXFovNG6LI2Mq4HkfXn/3lVIK/ydwVPJt7+3Qr1dXkq6YcvIZS
p8uC2dumxr18TqHL6UhO2jVCMYBz1XSyGX6+g6u53h/THv4+WjL0HKXQeD+xpo+yR8BPena6Arg9
v8BysvoZ5wXwMSmK/xxTAEn3zrPEWhcwSPCdf+Ecfs61KQ95qLvZVrDwAYyD98ZfXzTQEsnMZRws
oVMGf+y7W8w5fXC1stxabQ+5M/KrAtl4V7QgxbaZxz6f0UIvo4hpoPcfGohnwNmds4/AvNrJT6Bp
jowKuVJCAoK+TsrRaZIhRaH9MuTfOwn35ZsBxUlGA5rCHwy/kCFQKLUQswTaYnL2ZHrSbwhFcQz1
b+3rrZSoG/2A/D3Xeii1mg/NYeG4jzJ3y6+S2L8Rwc4CZl/px1qobsJfm65df9zqiGFZ767AiCpI
6dNApOMxXrX18k7jiNkr7ie2vGKEJpgYNfWBH+gUawb7ZDdDXrIe3EcXnIcbwN5JsnS7Gp+EQGW0
rtYQyOtytEWI9sTWT2fQkR+lpGt47KIN4/6Ep2TexXXHJE5jiI6Gv+5Y0UGiU0xNi4odrdFHWBYM
KRiKgACbznRFSbdXT/X/FSoGi4qd6SKY3eH0km7SLmSda1eVCSoAESyhZM8C7ERW+UJjCC3H1dCy
m7m2GFHRYNUR+SvYNRFIPIc64N/GoTpwoQ5gKqCPV/ZpF46YfB5wacosH+rzjrf5fO/1iMBHPa3P
yqCiuhR+7tSRgl8GCzgPto2j32188ZKJUBtsMgXj/49fp3JO2yBX4PyDf0rF0nm+J2Il7CFhrH+w
FiFdPLH/lfgZCpKZcOtGg17e3QxaY3nlRDnGB4tONCDOM2eXImQkbykRfIW7lFluVZwsxosjXdOg
EF21yw9LzqrXZsv558ItzXT7ZVeoHk6BPvJHfxDh/nd25L3AwfEr93wm1/Qj6ikKHeEBa+F47HLc
zegZfmpkDH113/EGPKXTlpVfylr4GrcxWoQpTQVS2qvmrZ4tn5zP8W8yi1pcd55G0ENxh+Qwvhqj
noA4dax792P/YJDIAKpI254ndRgoMSjm4azEkno9Wjl7wtcqs9AieqiFiguqlMK07FKMiSPcB20w
6L7ECbtavq1mIvdLU1MAsGuBrqQVpwrorKiWM6VwjEpd4qjhKFJKgkW+RG9DGakBz4c7B9Oq/nbE
3motRxj+0/t+h0jflWe2VMp0HWh28SkpXI+EB/qQGnkKn1k7TgjHT1blApUMd2mGlC0TYhba/dxl
i2GBFdScQPtdY1bkYPZpqGuOjxbtN6aml/ixcwKkOL4ck4YcIO+NriubEzKYjbvp0bL2sa5D+x6o
W9ZlSCP/8ye5rMDEKCsmG+oipP8QMViqFrRLK0Pomg8haB0J9YlK8OxCCfPULBWyMYWc6X1Pva6j
6XeA1GYiXbxDchr6WcnCcLaEAbRnTAd6BPanDom1MsZyvnssKTmRrgv72b0pAV1CR8emAM0tVgAs
XvQy6IjmxJhKc4cfEISF32X48uphDz/57QPTWbZX9KL6j5Yr2WBV+T3iApf9xXWBTIbAdWUoDZJO
3uECg2Gz7Qr1J5z9owQfeDDaFg1dsLNVpn2hiWXzKlE/FW4mUGX2JWaa5z3L4U6QkJluddcexIsw
sSdrLo4KPwbU6IH4hZ+xUzWI7xtbbNZGa2sG1KCEpzKcbxH4lN5tBzMYRppb/VkeZ2Q/sTx+abrp
muBwgg6H9NwvxI1coLYaFCNGN7KnZYIuXvkBdpj2B5g81YoMw8y7bpVo2UHH8j8Yeqz6L24t+Ccs
WIH894Ckq0vJzqKiERvf57J3NN317DoGWMbx/x8W1NWQ9IoC6bs06Q+DcrYVZGw6R5Fm32MpfeJe
B9gsEnj7YbMl7H+YqraFQi0qyiiZj90zYHsIO/96O8Uo0G88M3xMuD0tKgC/VzkZxL4iN7tL0ydI
46DnCcmkgJsJZuK4D1/ur43yBiSMfXnIlPY/XXZyyUzsYGYMcsOZjTmxRxvBm9eGlUwaza2TVfHt
TO6Yg3sHwiafbi/+mlH5Qa2gnnsrbkPslAPs+nDFmVWWS7qo2ufkdkzYsbxMlC5i9DS6lMf+LTJO
c+4kuwEBuRJT0NqJHHSZ2g427Z9OGm2LrZgCkRBPK53IEu5UbCf/ifEFt2EUlwPNgOL48kOW4ZOt
upEEg7KNQ2+RS3WltKW+5FjMbICUqHF5TX4JKhkk6eQiGPvpMsgMJR7YFqqO1wMw6Toc9sB/fpaw
Y3cnXF+yTuFkrn+Vue1VE57TVBQoyn5kgyEgU3IYyvZQGl/lqJ0F/zopGEEZ7D5dV0bEOyJ1VUFq
Or5TdJhDTTugxQ8NqybFqAmvVD7sqH7WKzvj+s8KH5YCBrfxkxP5KA9claKiGuSbk234OqHKRPCT
NzctpE+tPVXkH6cDsZJs5AEr8g8k9ZhOUDkADLTTs+eB//FzJBITru3GSmnHn+w63+wOfBO7rCMo
Pckd4ztOcud+Sol1KAXIVJvsPwBRq5iHTzyoZJvNiULTo77uUydZGNlHuca6y19lzyDSxbRk4vdh
YrgIZuu8jMHuNcMbU/lz1caog2XmIuU2EdQn513/mUu6YNZVRGzcITuh1U6yvbCfRmjQLypxNz6L
GnZejESL5GNAK3GNmHj/W1ZLMFlNdj46BsXJz1Mwo54Q8qigtJEoWNs+nv96G1JCTtQTNhcyGIhN
rO6PE+LT21DOFiai0eKkAGxONPliaAPaD6gGMe56cmmAOHpn3ouEVcqJew/WUkE624DTx9oyzzn1
zxDUmr+rHBlYaQyW6cHH8BMqmOCxg8y6J2yBA/mbqtpzcBIiC5C7v+BLjdPf+Dhc0FIggi6YDKSt
fH1kxU9s5ptVdphG4vBqGCnordn2vLg50ftmoPE+wH1vkgw23Cv0ntlxIB55x1ZTz3VK8gL4LUfZ
Kkmzcwk4EiNXCElAu/oInR6sTUCYIZKgmGW1kuld10uM3p4GKDfErfxcFKS7Jjm7M3awe3WmCjiV
qnG8VyY3QIIec946rmL7glBr/mgsZeB6jzkT+5z+7YMiTi7lFEIJhg75oBDSRaGZhljh/kE69HjN
QSAGb+60oRQXCCEKDid6y06Up7aWaeKdBg7ZcrqEFBc/pFJ6aznZuBIvfXb1J4zRvlx5GhqHk8kz
M3lwaTtT/gT1T4CgNI4heMOMNM4Olak4bDFnGwTp/Co0A5w1IesH6RzJY/32HHqWpsY3QjztmdxB
Jq0axsdLAjlQzfWEkz26NeF68CW4kS0j9rTjQtkUK8obbjmxXuiVURRrlMOR4OA4qrqLjRVLaThD
sLbRVnMK9ya9GECeTqs95RFcg9h1zVV5raVrZZP3ZyfxabyHSuhrdgWcxEmgTsQRPlHsj7porXZo
kaGesPPm8HowLQ0HMyXVbz+NwaxIUemsMWFv7RmTPOhr4hLd/5rh4//xDMVX1zJ8SWZy+YgPYbgP
rEs9XW+3i0mMH7beCTd/2slnhpPcGzXANSLrnalekQj2hYxtWNMm+r0Nh6uKLIqjMlZZomJW2pCt
BMgr09B40kE59QXomIk5szueoQ4TpedCUC+Jz1xonX4eVCEnen0rwahtkOcL+HhyqU9KYEaPALwa
0G0dpHGIjzvLENs5eO2opGGqxABqlYKpQtMh+LuFe9ULQWkELR1wdoKDUPlyfMeMUwVbaODizHsU
Sg1+CGhdWU7jdlmGMfaBNqumqFUImaquo08aPxUl16vfjGt1Iyen+hSRS9btYuGCxudKDgCNNuOq
Z56UBH8u2h1IH0Ecgsko+i5YCcrDqXccDeCJdmly+4wYoOZFWTC+gFK6FY36aL/X70TTT9zIkTp9
jaDm9Ox94T9Oe9RrkVumWTp9evRCVDcj5L+rhr6mphJMR4I1yvJ8SZhA4eYxI3AP5kPv5+Qz62bb
ayD/eeNxbRx5n4Q0GrpmpjpaQlvinIqM2yMQNK9AMJd2H4CYz6JI1sn5OA6WmBTHD8TWr7Iak1qZ
zhZI5jdkviLpn581/kbRFYwnRqY2XzkVTE22NVLXSNk8N47h0mGO8Gyhdieoai+Mr/XN+i0SrQIx
CO5eq7GjcBT1a07bdcSMoFyrPZnJYkGvDsYX/e2XNFRRJRctN4cWxhVH1GcROTrMGolf/HB+rLKS
XEBgTOnS9sp6ZpVe17Cvf97WJwv9WolriUQC9JZjoBuFitkq7l1c+ETeuqhuYFqxMX41t3TtgTDp
94lu4d/qRBNbuzwD9YOB+cHDJ6BxGshipjH3CYsnYf3+bwwe29u+bTfGLYPRqTLMb78LhxpEx+Uo
IC5mv1zMdASH/8cnWFsWo1lLfdlep6lOkkboZCa7OTLV1tCGaMSspWR4c4glGX34J4mbLQrBkiRn
wZ4LOZfEiti3e4xXa9E1W5fVqp2Lh7gxosVcPpLiqaFvut+5B2vHpSM3XcU4bksA2doEN8q/B0qN
7+D+tnFxHD88BxWEzp0Ln5gAx58LeJ63aWO0Xk8+PLpU30QW53P1rfYYXbf+HfYiqssS/LMoPYVJ
rbfiWrC0aneVdmWSqekYZ4TkNwuRlZyx4sC/UJDDZHV74KhwUXilzHbGataFKvgsdQ5wkNoAFIUi
B8+9QM5Rl0QdBBesCzChSjqmdAvpUY+XRWuVGHsfJMllcagzTA6AGhz8rfAvI0o5h2bW4Pc34YuR
9RPOH1uXf06LJLT7uGOhZGxMasTnqsAqDCRddyRfN0efTfIA54OTxauUzhTyiIYoJ/cnBGUIHO/X
uwJdg+cG581JpVK3S3moQymRlZOBqTolZlXIY6hFYqZzxrUvjcdDuwZoHg9vVoK3e4rjPz4IeyAe
8GOsjvhiFMfJ3cgFywBBMmOHTy0ORMtoCFnAHcEgI6vSYSb8z6ju0F9xqgftHEt5POPu3EbRmqmc
Jt2FG4HqKhJgQbasn/80Wruz0XGGNhM6w5+wROSW5mMH4HrLk50sqoNR8/o9ZOZfeUJTLDnXCEXE
c6iUIu8lFg3RKrhKhRSH1Ne4rDVRAGvAX1LF9vflD9JqIP7HCMXtFJNOEwKJk1T8Eb+uVFCXd05I
83FOsrjg8p+YLoa7qwdyEvhHKUhHNNZMOauvxeYT5JWZlRb7R60/NdsxzfLVcd4XWrwyZJDK+78J
G/AEzQ7BzC4hppUyyln9TLZeaNt+SKGbHKRwZmXKU97KveOcO4yXSoG9gMdiFqmE2IIC84uFEdHb
Fa5sMI7meFI/37KE3AHwxtYTUS+z3Z66HJlnssrZ6Uha7m5zTWv8HhaQO56r9UsTfNuNjvvPaZR3
UZpOz8wM0E+4wrbqnqO9y2PFwamC00bSFlQBiTnkTLz7AgvYPJuRo9QRKHW9Rchk9+MdJJbpQk41
BD34y7j92QW7/kxlakLb2c3jjCGgv+26FdpfhRTqYdnlDNv+swWWmNJviyF32tEqQweWAq/c3F29
K50FJTwycEWqPX2dcFVvXN1DxT8hTzaESEOrL5CDHCU/OFjP7M4+Gxj07vO1L0z+BXibjMmA25Nm
+N5eKXAh1ANIpyo7tQw6UI/kamWxkdGCPj9rZGhP3wMHz547rKuq9UbbSYN6hEdO/1aT0V900F8e
mZxu4ROMUp17syy88zMJ+d2NODEw9FrCSU+PYzdI1D+zi/9Oqs5KdYT23wchp0PgXvlBBp1/UaMG
VQIYX3wyNLAM4KcgJbFdThh56HgWFVnMI/Ae3ytuc0eRhYMhaGiGY/O9q0sL0IXR2tBtmAyCO07G
xtmFyaQlmLlCeV2yJhSsqxA1tANcrlZhq3Xf20WsxiDlz0475a/ODtz8z/uANm9HATvfviYEA4xM
K9l8/+9p810iaR2sFGZCDSkpazQ9wKxUuyx/7p+roMMwjTPqhFgV8KdYuPznqlIbwsW1XCNFx0Cz
uzhQMoLw5uDbuwAOnhkSi168do0nigOWjPHmpWdvQsQv41HBQw4qj/sQ7nw1phkLZSkc4vev8HMO
+hBceaslHnLXGNGxXZNK7yD3JamA8fJ1nQbtmpqugINu2hrIkrTfArFTs6+RxZaeYnTgBis0YZxN
Gl05qiNeBLuFc2O1docCJY7YRvnY31BOXfUtzyx/24FgooIzei6//Zw8MyDeVSETh0GoJ0zntn7w
4pU7/01DQ7nV618IdkLa/tyJsGo9NmkCgxjqw/99xlII14Uj/ZJ8oYVTACQbwIppDE7MU6kRF+Zv
XPcoOI5z17xV4vlfmC0WTMbLUpsQE7E3n63mSnMBmYliX5BhtDlOlLZS7MAGSpPnN729z/IYPmJK
FcP0kKekSXit0gXyv+Bxmd8F7Zw3g4OH7W21NyqYPVBlkftq9QZTmDSc0qdSZWwXERBtbE71LOCQ
Y1q4aUj+FetcEKqDV9UJ7+QWGq2CdStr04H4mlYJIBp60jSuDa3AI6z4OZSueLnocY794QVtNabL
kKmZqNUv51m9T1qXhw1D78OfpcUgctbNPg/sWuzItozx2MHzMI+Pf2v75j5mqC4DwBb6oeHoGBv8
iFLgA8+YFSNM7VO66DuMCD6U1DkLlb2Vnp3FzcgLoqfCUOZkd2QQZxSi5wnw5sk5RU21ZNfu180b
hd2tbohu30iy8pSh+S6UkAmPGoLIK8dVyrzPG+tiMLA77MW/2iTJzce94nqwmRbnwwz+1xCG3XjA
LpeN2XEIDzU1GSAgukATPD3kvwpCcnpRqHBQpZDiEzcwWRMTAqyTTDS2E/3FGzxcKcsDHrqypCFT
OeTCu5qQvaBC39RO8iXBumPPqSKjNDPheRfGD2lIASq8RPmJ+7cAoyTAQox4dl7fPKfcJw5q/7Ij
2sG/PhNqVnvzVxVn1NwIfgCa2i+vOrc5zQM1l7Dp67ijYLJPX2YSRy1GyPCchBMouwsShdfbZM/t
oSCU1QrLKW5dxQTj+JTdCZYS8GawLsFDy4WIgWbQ70Dnxg6hB6Eh0ou7Hhe73kiOQwkhoydnBeC1
KCNHK1nupnqkMNZHNKrOdOg/vM2Wd4HUB9PMBmXsu+M+veDuwpdqqjFQfIBR1uaCy3vxZZCfJy+C
hfCvthshDGPSTMNxyLzFaXcKxVSuB9APyLzcp9JnCvjsjPRtFaHiNeKr5dcyhloPFc6lfoDiecuC
ZLP3Qf1xAXbuz6xXY3cTr0kt0UY5Ed/uREfiTDY6r9k7GFx0pYxmxroUdWVQfWdhH3B34LHQOlPc
uL6NelQ2uk0VE0sRu1K3DctWwsFjQ2U4lplYK8M2MeGc4RLpOLjbcE+PCrTWa8CMovfEOKCstX5w
6FQ8ddmqlHQVl9jXGU9fGkhfSnE8Lx5HLjnoLq6An0OhpKBNMiG8JB2x6KtMQKMo6+//4u9+Bd74
YzQCT4/YG9F92blMu8ZL2RDT+nlD9Vsbkzdkc8oC0ifKih0EZZi3gjrPuyq3oIy+42noVTCP7Zon
npdXQBFyWekrw3yWEFW3Slh2qtKizju416ds1r1E5vYrt/IpVc5ryG3vYJXodXGsnCMxBCekN7Ks
Vmyt+CqSzkbOZO10YQPafCEG5/N233oXsB+gWrasQO/r0i+6fWo+deL1vCJ9hJkW1934HPOL3h/l
/hGg1EFcgPe0K077UhDExl4Mg55+tfyhDQ+wNRc1Krc5Pfh2xpN8v03BDgduqi1a4bhYOSZKaP2c
zljvL6iG7E3ZzLLcu+PzbI8hoYXAKpSV0IIQgM7FECCbP7u3AOV1TO0ou+br9Z9LjBSIubn0aMWp
MIp8MiqGzjBEbWU6QWLBqSuabhdDgiqc4nHVLEh/Zs/5dtxIWZxFQBFHciqZoI5K6JYI9DXK+osn
svW1Jhpre7pPJlmZYSO1pSmqzPF8V3PfrJHwlfjIymUYr0P10hdIAv3wSt8VgSCJLOV7RtflyS58
elABb61n7heKfLdBP+XdU2eKsEjMwIDnf0Mz51HOFTCIsVtvyRHKNR+NcNDgoIy/jZ3oqhmczTJK
u33rRrM7QTPkjtyV1yoIiuAeS1S+Z7dpR9UTFXZE9OdGb+EDPYSL9b0iWi9vj5/OpdpR1zbF47kn
blhzccCVakGQPxTRSGy7s9wo3IpAAR8yEmEOksLGAjrwarUQHcAMsQvNAw0d5+6z4f8k2XgRs1x6
KPncHp/26E7OlwBQgEpFCSoqHY6XjX83186LYWuladD3whZgtjRRN8zK4GD8bdSvdIbgxv2eV52g
rKz8QAxh1LrbfsLfmK4SRXWZsDQ0FCzn82c9cEynoitQBCr7UwS6ZzaRAyLwElTGfjQhdpKty7os
TSKBmiEc4dGwCYtalsSrngsA3e4N89JYmcZfZ2IPT3PvsM7JMQ+J6ZLWVd2Ntccox/WDq/g2S6m/
EAwz+x92KVlqeEOalRWYntGMuUMBCmhEUjG6XBWmMb83WjfSXJUQliwIo6CAc1qhG/mhuh8w4eyp
lpYRZDWmMJ3/l+djcngXnGhff+1AeMAHHFYIRr0HZhLydex0FMQ8ZEnTmP5FAx9nfpy1A3YnJJc3
da6qCk5sNBr3J96z8JSa708eyrtjsXUlBwvsOFAGPJqRJub+RhcRNzMQkUaeyxVk9uTtIKXaQgBn
eTpobO4baRbCt85pbtyw0ge/MxMf/OUClMAKqW2up7wQWpOBalMq7matd/utN72f/VWluau943o6
x9etQ8RY1DJwEQbhlHCaL3oAOqixtVSB4y7hK1SOOIjWQkD6clLzAIqb//oQV8RqOs6qCzG2YTzk
zBIw6C/CSV7Xp5kMi4d8i6BC90jn6pjuI691qZz3PBS8sE9tVCBeyCW5ZA9SEUFp5RYEhGwPidu4
4nCCz5EwCFvpAq30sVqoR5LNxsRC9bdAXlknwI4E7MN7iMeOrvB77kMPVEXTcIIffCHRkUzjgtoT
9gq2O1rQh15uH2s5I4Lg+x+Oo31slHiqt4YRNEdp1YHAkKzlS4OUQMqg/m4V/PXEoG9F9Xkehgv1
w4OfSv95naHb/gHcmL960X18W1yMFw6xv2v+KNF0QglAbt6x2xBplwVFVbJemcAAE7BlAr3xjB1U
Pjuo/+SYC/xVa4as/xFOzg3nBgvLTK6f6KpA7s7Gudy63jaq5o7Z0G+luQEh1K9uz9wbcUkilU/d
uMPH9rCM2Neb5MBsjw03t+JAdQkdsBraEgeTnxLIt+pnx/MFmvPNf6LYSSeVod0Vlks9uSFNqV1F
Lxzl7utOHwyLdW3ZOdIjLpm1yZF5TpyoDceLcxoBn9JGekYzA0Hdfi0sLux0Na7XcK8rMtXTHTiY
r+AaUduZsX+VPtjkBcVbwXqagVu4+jRKLPfudyo4cUYSfU+kusYZJfYxeBMo/yXdHJA9vsBHHqYS
tB34GtrNFtcudwPIOnrlolLvSQOaOpdX2cs1+GDXpLVl6VJLroToh28wfDIQtbovIH5bs7Mov2T2
cumBp13JkvC5zifFhHvtumnkbAZZl/KtAQmOntxcElZ7AoGL4GIIgWpfOJGkdSLnw4o/rsxvq/di
7jdI6fP3G5ESadjhVeN3Vd68HatHIQyT2nIYUOxMZs+gD8z1YPcBFAzTQlGSZqcMnLYlB12cCiQK
3UDojmAqnESvZFxwx+g1aC8fV9cmEroGUO/YqYfasqxcO5LVEnl0gwDpVlDcDFfua5eI5MAfMFmt
+uyilJfYUgQB/QBHtVNvUV55gmqqU3coB5jgZ4K42jmuVZclPwWyFzfF7wy+jvXqBs1jrFKxn9gj
r8TINyln3XOAL2v5jAIRLf6H96ACMFlUzt80ZFeY7rpcp0v2bbifQCcyXWUSB/TnJNvNfLd8bQg8
TjX64HyZLRjMBfWMIYSTrkCTmABMyDuhfUzEHvKZFDWNP7KiKxko99nn0lOE1qfoyZVNthKIMK7o
ZFI6mEv7zINP1jRxbaZS330Gk1q1tTemma8z456thakPRFAVf92A9XusTti4OGL200o4VGW4LLmP
64dorfx0AabDBLr7lIdtl092iNhYIyIqKyjFY2W3SIxozQthdb++Ww7NCa5NWaVSRJaJMiz310rt
FKqTlujuE5iBLNaJOM7c0ShhtUzW7iWEYwhtKSo9oNPSf4WnburwhD8P07/JBtmLcuyYGaKWhqv/
pXDCy72lU/eJ/u+hWliNtb4y2IHyYkd8ce12Ie4lgPp7cvPHFtHSJpw7kDlK3Sm1vIFVvDxf3XzJ
uLebdbPx1m9pXWknhflvF98IKG83CIqmfOshJ9kkbasftdTVJNZu05XdbNBnhJ0wwt7jksQgAGNu
uaCwQya6J5r2XFrc+Jvhi9eJ/N7EOEBDQYdIDOVOaNWkn+eiH2UYqgOXfksv8gc57oGmhDg5AX0B
BNl0K5ra6EpY89x+wlxu3CnBucAADtKaIahIKgQ+a2FZQUuko08U4FygOwDPiDbbMWTpvxSz3vtf
kGu9XCEFLAtJRHvvLntB2n6D6UJro40zFjjYlDzskODp2xY1gDCsHgtJDjg71OnRzsTf05zJT8Oo
8Jv2NDe7kQQHGuOotQGpABQZpe4FYo6MeoMwSbq6R1YDj/LWwmdQeOX1ZTJ9bgjl6FIMmIoVeUso
CRnwFTNEbBN46KwhxvDl2D9p7U3Gp+xw0o0fSKLW67pqgbp+rpBrJW8lXlZodIBjwXAzff8Ng13k
hMPkOn2VOePTR9dvAGlvF0yC1dOcmM+3UG7bh9KvZrV1JtSIYb8Sk5ox1V4rTw70+KgCAeMNqGZg
SBe5uuuCdq+0yMLMGb96zsSY1xyMfOIbr9jlnUrZIJHIWfHFyQ+lSNS3q/DVPVtepcdFcSh9qMoO
uacpRlFXz2gFW5tcCNjPvAWKmTjT5Bp87UWpik1foyvS2H/62L1mLZGAbcya2XX5EjCG7l27GANT
f7097BZgEVYoslofiR3KdOEZpYBFCxA/QkgBqI6LLRAvAelMZjhJ+TA/lyvy5IpMmNDvf3LqGI5Y
8xfRKYWdqeyTwIxJkODv7PM00rcQrWwEELqC1hlz/yCYkZBc9jNCiQU0lr3YGfxS+g+3C21c+Wkj
/8kpbBvbaZBHDzA9p7/pDruPP155OEnfiw48TVSTFxRINjvfHmCg5O0FlsIIrATI18Ov99/xr/q2
sDSqUMqPnjckYxsBYSfhbeTsKLJEVMe4grlMUufa2NXWthjbOgN0AItZyefksgUA/ha6IKKyVqyP
/6glIGA7M5fX5PNx3KLciQNtmfAd/wcwLeirgWW8FrlR/l/plHdHMw9PWt6/+59yjAC9S7m2/GIN
RkjA0udQoJ8cRp+fBzfsP6BJgY5JoVynBoF1XQL1beSnwXOP8FY/m1yOLW5JMp0B7Tmci3S5uigP
sppe694bMoj8ci1wU2+GHGldJwBmBO9uz5LV1DqHrtBA+c30znw/Z9nYUdkE3iQw6TengOtdtfCB
NRnWCHdjvOcvD+h7sDhHfxvYhgsFaTl4JntElziSphZ698qb40/kzOtqoRoE7OGknzW+DUPpj1B6
cq51kNsbBmeB21DOQKenSJ5RODxGml79Ozv0Pme1moUrSIjqVjKMkZb3lRpDBwgQgBcuhVh3lgjB
MM0EwiVZK8OSH6jtkgRPlPxZxpQl3Zcqv4F9LWmYJ4KA3+HroXpGnngWIRNuHyTvJB0PW5OKZT7h
O+OuewYjHlWabDNpgsrBehwScxlc1R9m5BPaDhs3POBmy9hklTK83J+sMmEsR/fo4uT6ux+IqjSh
yUlhdbBz5GXDYR9jk45pJ7EFn6nDddS87w+cWYcQFgtOh+FRaPoZ3jLSeoNepfjpnsim0594AiIk
bgA0TXkFXOOG0d8hD7LTGnJx8B8xrENU+kOHpx/AsxzlttrxUiFbOEP0LLJfQYOZ5nNSOf1fHePx
clbs7qh5fP7vOE4ORRUCsFFm+MByyTYFkwG6K4RaQ+SA6In0yuGcp6S8Zz8UnmmNZxJTtU6qg0D4
Cvhd++i9qQoYceLZ1iVkGmEbYuCbtOC5HzaCpDsGvDgrGCLx/UO4jpaf6z6KF+i//FBjRFIQemfW
KCfFz8fI5yVZwQsZSM5CW2hlZdRhLtL0YPEE4b7eKKmPF21S5ys2E3jKE6uaibYQSL/4AX17duAJ
6klOf9lkD7SfwlxE9UBZzsyOHlBZ5QHRlA2gp0ELL9UcFwfBpqwfmkZbOK/WcRjTxTTZR0qfvjmA
gV2JO3mE8V3FLyROKz2GvXem6Mp7/Z6c+FD4L9wAJUmFg0blSpkwMWi6XSUym5WVjr5TNwKEUAVw
r5nPZJ82Ot66vscwc8hw/lnZeYkBZL9G59URKkuCZJhC/FImUzyhCh+Kzfj7k3/G06VeRWM/YLdH
oA4YniGz1UoOhehRSKwq1qzl74Y9qsaY8UKbacwKS8xiO14PYO5BHxg6lWoAkBa3Fts5snGxRTB5
bzFvfTe+uu+HkbtwZnmWHcEHlc7I0aKdl/vXAsAaogNYPmgthItdu7l9gxexlnJlLLZQnaeLjaUs
JEIF8+y7FxjHaLm/FMbHkyXxz3ZXrDtFXcbTi4SR7pKL1hwuK9AWNz8POXX5JKUNxLNA6yU0UGRr
oZ1ZcFs+BhYbthoosMrB46aU/3zIopfUipcUWHTUtUJ9B3PF62GNBVvMfp/4JK+WszL5O9BkLhkd
BZx/2/T0SVua+IiMIF/owks1ueApujrH+V+LXNBOpv+5S+ul2YrLbvYxCqZlVjdu5vzOACgpDRHQ
LlXZRfZi9ohubZlkgjx5dAqKcqXkLePO7YA8tMyIJsCWvIO2ZIH+uY+6Q6WTuGsAdluPlF+GaIAb
MGjARErWcdsdW5E/di+ugEpymAMcbWYjikkM6XTCQfvRxCRjGYhzf2aELdyzCIlu9yqyzFWrv+lJ
ZCPmEpPbk65yXyaA/ZzioS8H8wxWQj4n28QNlcz1tOBcRCYiOZYa7kxjVE1/Awe8saF5gwOQBh2d
XgvF7KTd7axJL+v48UteQZMbmU285r8Br3EGXDRp/vVC2f9f5crgg/J3Nw7/ow8Vx/qs0YU8zMxl
0bdei4TsiMc92Q7ujYAacOsy5AxET7OHxa3YzYOXdJah7/zd757is0mOv2pU/fKZm5Na5PVoOwxc
H9IS1wcaWKYFIVkHyvWrMu77uYFv9AUCOYCl6PQXMaz7gklY8lnAGP4HApEz0SBXbRnhYDdQ3Yxq
s+H/azjgOZSvyxak7t3Q20eKi8gE2U29W5eEvK1kG9u/AHWyLtD38Z5MrqmyBDZawrf8HnlC3wFr
AEH8yrTBmf63TK1oh8f2Y+lySYY+2y2T5ns7JISD74JCLuopSJ7BjjPgPGIe8lPrwh8+Fssx5NA5
PIzCcGXDzGkB6p5ji05HAXD3JCPcNOaB5m7kG3CEF3gA9rR31X2SzDjw8IPk6kwIoS7goMhIqgUs
MrStoj9NdXCq5ErH8/OCmASho/McKBdIIsmepcb55NqjO9z26+DppsNkQwRuh0fCkkF7Io6rl8we
tv+fNmpAVeuJq8dM/fJy0CBaXsDuFnbUtavhVyNsM1Oky46ig3rya5BHYWfPlkXJIgqdHz+dPN8Y
/RXF4B+33zcYDi1lgt/t0wSymgAWADQi9WUqNIbuKxF7gXD4Snq02Vs1+xPLjzxmQu2020SdaU9q
yC22glnoT20kFxlx0bQTKjG8SmCLSunWeLI6ztoSbRz3X2V0NlEpYAPyyFxKo5KxOAvUFlef0WP4
NXMR1XxbnhBJSi5gpzlUb3dAzW1tKwLtCa12qLkE6a9FeIh/ShIGua8vt915t7LyrQlb0BR3wwyY
/M3TZ1OrPoQWRTgLsYfzGdyQdVTtuEFvOU7t6HjC/RwXI1HlHXZ8JpMXTu8eTbNRT8tF+7WpsZCV
mFbnGi6iAnu+pivKKCNi4hdPe+XD3n+IHMZThqv1yQqjby8Toas/w7ZknssD+ntrGOza8gI1oAc/
08iq53mEKc2/RFtog2wIj8txxuiJifb2etRKNuNdm3dWcD679dYdJwWGzCTsx0DM6C+3rkATV2jB
lLxcEZt9kg+J9xW8XJDzgJT5rtW1Iqm+9PY/4K+xwg9hqgAtSIMoWJvZYWgLzjlmZotHbfixvao2
OgvHZZ4Hv6oVl5L6xS75L789JXdWT1KTC4JqewCAusgQiUI+2OMEKNW131vmraqAEvIcHNATA3Wr
iafiVb9Abx0oF6iz7S8Gx5SaIg6ngYN5i9dLZtIyJgvr2WFaRsHvbRsxHEdJ7BurdSsHStWw7fIk
zRjhZSP3AJv9iVnrRWSspNO7TPFGTXlD0x+Lhk2VNyif3yn1InQ/UlAp0yB8gVMjQDj5Q3rnj3WO
Z8mWGCM460TJjCs4uS4n0P+kW89f5lm0m7wIOgPd+DGekioXZTC63ji6WvIkVZTRz664IGmBufmk
8vCrON2jCoYdVD6VfEzRlpE/BQ13ETAOSWJeRi1KBOSV995y4qyODdaymY6ZtCiFBU1kzJsTUPCn
xL+gB+0Pr0JOaME06D4bLVfB9mvPtnDgX16VG0cnq5aA3sJpexAmaO1CzYw5jqaWJS/Pbdw+Ttpq
H9OkyuC8glLIAUWMn9q8lnSp6cPBuh3qJ0bdsZ6vPjgTynJzEJ+33UaHbiUqT0aAzcYQwaHSJ75B
1SV9IPSU1iriCqCtUre1J4WxzLJCptMjkTdBfzqPQ5i0oguCXd/DB4zeIkuWY4pQXhh7fgPoxHLf
KI2lgTtt454AWzQ5uIBZ6/xFDOgnYQHXlzoJWqG90KEzzU2Aanpy1AABvRE4hZwPDPifUk0KVyjh
8hK/9im2De1ZrF+QxiEFyaqmtJPNYWFiCPRnmr2sFHBFZzQ/dCd49d+qUSi4POVBPhXQhZi4iTBX
sElniBxC81rMqKneFdk3vLH73Sybx7A6tUCBwy2AzahuucthXvaWv8SsQVUdQ0BRz575VuWrERwQ
FcypSvGIroJplKcAWpVnlwuoxTm6ZPmeXDFjB25QB2AZku3MqagYEHlLOoTy3YPoloLORzxOyY6R
zoT/aU/3PixJaGHcGAMQtL/bOV68fWJ/AUrrXH/f6w8sobo7Zr2XHkvKvlMOK+OCsa63oP08blJB
Vr2Au8U7LH6NL4dW23+50OcGbWrmOVDK0HObX8gMjTBv/vl6L0qCNCnSIIzT6z/6a1gjlyHrqteX
vOZWQSidkUXZL1CJt+xv2WBcOooToGC7iGW6khwhgRvOElKUBJRkrhGcmhx6qdxzK2Xg1Mr6ULht
UfanSTU1V+on9c2QhOK859Co+C1w+OJwZc2OVziCu5mvpIWsLSgjMScdqseOJT3X/hQCJr81IjWN
1IzpqTwgfcgE0UHIxfQbucvong56VAHfC4AJTd0AvHVvPYVTuHDt5hd7U8f6hGfiurxk3zFW2jwV
qe0HWl6Xiugc5MARGed7iazvC621h4jU1Nhon4SCEUVK6PiP5lSE9iTICIysMnTsHT3Njq83cT0L
t7xPADYinf/Xbo8+pb3R3e6ZHzqrtVFgs3dV750fTp6kKESfREEz4eUd8gcIkFnsPLu4jnvtmdyI
0m8Cs61OvSsuLIAWqMk5reP7o9Ke/ZFPzkDzKcLAXIlWyr6Bng3R7aa4IOQxDmsJ0uC8ecvUdgnN
9QD6Wm6f6MzCWFBakiK24Rw7zL8WVIi/EVZ5yYaNC3SaOzVpfHTgknuOQC/n6h/75PVTCq9sdqYT
8CfV7PdUM1OeGJiLgVKZcindcpc2xwYutvkNfDnoTqybTwfd9J4u0tD8/UyZCPPn2oNFtCEaYQly
CZRhpW8TBglyYd5XIwnGQVMOPHD5RwhS8gqVFqmwXwsKNnRyD+DnUhjqTzi3JEY+LVHxyNu40335
boQ9viuAoGCeKFOyfNEWaaMPmuKiSICxxu2eFty8qn/c19AYs5cQF7nRl3Grz07YI1IU3Cw2/gB2
gdzlcHv6mit6ocx9Tk1Iz3CVOAxMdZptmoDqsbiUv7xaiuvZviGRDLTIXLmOu6f9kB6wu3K4KuII
nhbFcPdTBypEH6QARKeTKwMN/8/eJO2CtlRnEhHTZ83NtRiBHTIB8OZvQuvbuMhUBfvg1r5fOjX/
CTiWdjTyyYRUfmiY/uqScyfOPHpsHd+Ylr+Z8gEHpTGbzk2/r4CeAS+fCyurN3jMQ+sfAxTPA8Ec
CRtxWcZE7rB+RQRi+dyQB1PA6Ynnggem7+BJuatUG0vUzsTwMuZcgnWdetIQkT+lu1f8op/nlRKg
aLo0Gqtpt4LfT3/H5sZw3x0pCHk1hr4TzloqmA21EjNflGxPK1lz9GzxHEzEFvbnU8qce/THxF6P
PFwKwngCxGWpxp6qee2INooxS21u/fsYjD8Fgz0HJf/wxw9hjatWp3ixB/QD1pRY0vU25+a9yq24
36QLoThxvJwGiZI6TZdubwdkTZPLHtWl9ShiEGAQrVpNf9hT1yea1i7/wXRetJYqPYE7ZiDkW3Zd
f1Hacqe0og25UPdwfqOgdz0EhNSyiFR0Kg7TwU+fOyCIk+9f0jRz5Ha93l0Vh2dWRxIpC9U5uug5
jIQQ6OKJBXHZ68PXh9knyenAF7PEd5DcyNz85jrFaVopg8UDbNpFcgaxpumxhdFk/OJq35luKZEE
D9jD2ELoeh5NTT7NpZRmBeWun8QQ0HfqAE9ei6+S+c3dtfZCnjKqCBmWBVU82gheNxuwnilHgzDW
as2DJB5uR6oHe8XRZ3hbg2exbziay28mWeVPDSAh8Y4z8ysoqWpewBhGuKuJ5nqkJ6YmiqNl3EQV
dsN2IqHjGw5D1F63EWT94krm3NI9hHmdxA3KgDksPdKzKnF4euDux0davLZEZVx2jKrQJC4SXcn0
rKHuLFrkThvzgf9JbSpH7FubFazBQCvnPQKkhvlfSm/2k9+mMmDkgEPyWEqGCdF1a/valbxgpyyi
fusAdyNEEIWeXY7ImLQm61He4Np8m7KijmsNCoK+IWDkSRcZlsTjBJOv7uThsLYoxDj0R2vMpF0F
LkxI/DvI8cRQaOHhuizFM9xATc7HdxlQlYJhufPWNd5XkzZwW7GfDv8ry/G1/fgI6+4raY+bqE44
XsIY/00+CpotWZqGuY1Q24JAXwuM6MrebR35gG2BdkSY84saSTfJuiz148TuUR6/A32fcGMjDE9k
EJx9KtJ9JN0o9M33iiA+Z0W7iB2R8ySqHEZs8mAVu8KYC781SV4afoCnHYRXdu9fHiCiQhn5csxV
KIaSZB0+yW4luPrkMFOr09PxsyEAgPI2B+WidqKTFUw1ud8klOzclcl/qN8cHPBMaIi7VOpjsXzJ
DwyyTT4/7e0HaK2FQtMT4MMkQ+hiCzlptkj2t/mSjBaEkmlV2H1+H7C93Cuh0NhnnLC11wsAuDnp
D6dGz8tVYbDtSnWvk/4EFe24IcTVM+SxSnYwKA40ojDPV5iLKbzBx+20DxlmLujwia7RV+3q+juH
5BcSWOJ/85MDmQZOhIMQJ9kwZB4pRT3CRbY2ePoSu4V9s8Er/oD+bzz5hmWqMxMF9r0FK165YDCf
Y2K/hQDGCFIO8VgX/14yw46Y1I7B7aGSO1ibblVRLChalWO4TkxmVeNQv4DAFGauSeNiCLPBsj3D
DCMnHtnpm4OxrKHI/xDXdvyhTtmCfBzSzrPH3+IJ1TsOzFdj7EuXZcwyN8emhOGIHBlLI7d/qddM
1Z8Q8k7nOj3xVIItudshsSEpVXjfhg6khbPLxDM/pwsWPacjklAnX2Uen1n1ER+ejx3FLUxfBjzA
FV1Kv9w3kSUIuwJnRq+H8rsMXMSzSOm8RBfm7roA+p0kCNDnR7+rSdPfF5yKOgJoANH4K1a6kFmy
Zr4ZFoqxzJMenLkKbevEmWAMLCfS4owh5RvIQrPaEJllLwB6cDK6+EDzWMb/fEsx+nX6ZFAOjo/w
OUr0h1E2wU9OD3VcpFuiB3ufiBWgZyrqCQh93ibIi8WVIW92uNs3lfhlb0HwxD7+Y8Q+rhp/YAhe
VsRd4BDQM4EnZZwG/J6s3q9CpYwl6hV/VRL4TEciRBPZYlAvQmlKDvdbYcazRs2D9CB0T0aTI9Bf
FiYxU0YysvLIRmBDeVWslXM1alQFjEvQn8sPSYxiRyIbACy1dKBHduNw0MSg8JQYe7SI6y3ewrIW
mFDuxd2bvorFH2lfdQfH7Yae2fNvy7MNjEbMaqp7xzqFIXTm6zNfhu+1CMdlw98wPtsWNlQuSk+h
PMY3j1312sKuwYqMKZWO2JCSqdWgJo0DfbaEtWfAVXS9nSwi3YgGRLkWdF0bGp305uX5lcxbQaXE
JQDKrawdLc0ZDbZL1MhCFytZs8ipMKAGhCGQiHQSavpwdbqaQSvQLgn098aaUSp7dKI2TPPwCQQx
yQJw1sJwFYuHb27mKT8L6ZGlX939JYqp+RXz4riPN1tibM//OdYc3vK1PS2IbdgivVHubOF6fwkU
jX5IJTT5YHbrKstIoI3ictGGHoS++4HE072KgK4+s+HHSr/2BD8elmoRJr7bUR8vmMuxhVty/Ie4
8A4XCxEDJg7eAJZ9/+mWXCc4xdnKsiP9Sp62jZBEmDUkSqES+hYq3ZzcQXk+ZvsEuR6OpsoNNKkQ
3QmOpIPbAv0t76Cd/XEqOMHZ1Q9VoW3imnkowuHFxnmdKrrDxEWrbLZHnySlb4a7x42CZOFm0uTw
0wYDz0tpODHCldP/G/wgXp4bEWW37WigJSmJ93apQZTV8kffwAJMjKdmeX+Iy9SyT3RlC9s1bdMG
keRK8THfrUXrzGUWN7CgNpHZHj8SzF97iKfnXrzlghkTI/Un1SkQDC8c8Y91i8kZqtlacLG7NP5Q
xibWkijMCCymCzQFNQ7hRIwLbgGQDBJEMcmxbcgcyOXmJfbj6dW42sL8taif4ouGEOwnEEq1SMiF
CyaeW5P4fPNX/ZA0hAWq1pnbdkJS0qkgOG0pK3c05flIkk9s838Mlz0hAz+KfxdMB2Ub1o/t72Jb
/FLJWnwIlEVl55Dyc07ob69T0p913z9QRuWU22SS+vWytqoYNRneyVBgXOhzjliIlY6wLWXmBnAo
KokFLLLfs8o971y1DopzNAeBo/F/mFqAT2BXw5hhf9mOhAXpTNcJF0XsKmq1fOGzNDeYKEcA5oMy
qGWbuvsZB37nZGYXOuNRiF42W/aQ0nd3Nu8+kN9ZbaNgsJai0uJB3SE0mU/sfl2S9SlfVQLHIoY9
Zvq18h6hDw/xjD/GFIJsL2FFyDjdajLeaDL4xWVrDFxonozp919LF0qP+ckSEPepv6GGAisEGfiV
cZEIDW3zVB69OFCfwj4BpzvFh+vvhCodWlx9cPY+O7ZDODUcwDs0k0lpnwl2HNbbOvipz14LQsda
u+ZMK7uNAlD3ZvoEMMa62nsliier5GsPF+v5Bh7fONdHgXk89H839eeUR82A2v4v1euXxdx/giAM
/zeDZZW3yFzLgUUsmS0t7JHFhIo5GTvK1DWXgWmozOooXycxSdFqrMYjHD8sMAfMEcbYf51VqZov
NetDpN7aDO2LvtqwDyFv3xljJVvhOXTEnc4Fk7IB9EFeitZNkWyVjNEpwgZK6eHiFWGta6dvk+X0
memzyunN2dw/BdiOCmuxZeBmmC/qFHBJqzGgzy3kNXOK7XGXGMNoRyiyPU8rXsTY/c8oMicitBrZ
SutfkML4oxhtmGqncvA/Rg/0XCNtHfK09mxz+LwH41JWrFxbNVYPdu/vSSYXvj54zk8IODHSyfjJ
9cv/p2zQ96XW4DZPeQm0Yl3V4sw11qE/iiW9xqQNYA3jXJlT0k+8/Dml2koZ+2OBynYjxmrUUFM/
yO4XHdaabopSPVulDV0FbnKcsnXareLTCTuAjL+iuG/q2DPLmC2kGL4l2BUyTm+5DCfEUi5+uxhe
IWLb6OI6Gu0hdjVrjblJI9+TlsPCnP5mpx6gpnP+aXAsTNE6+NWy/2rHElZJL8raXvGNMCDMAClh
xBVqkLaqLpE2QpknRVKFM7uI6yhcz0wciP4dwsi/4DQJU8mJe/zloRF6yQd8f8hBhzeFoLSlXxhX
uMjhZUGRx2TxvzZkTPqADp+ZqupW7pDM/XvGLASWsBdyY1/WwJlcuk0c2d6h0cFsI42a+7LoofQ0
rEgFITOMMuTqnjruwwdhvXxZCWVz0WvmixnrsDSqPcwY7MAKU+1o3zGG/I7+Xj4+5fiSpy97mme/
Q+gXuwmDQ7Uf3DsUJUE/Mj6EvziIBIwYFdhz12DHW176/AA0a0p2xR+TO07nEPkpREWRj24joCMS
sPKWbOyEHWULzBAu2e00VI26632hW+g7ot7gsXfVjrEfL7oVTYOzX9OExzv9rvifq7yNCNMIR1B+
qxIYGbqIJwjbGBGjPoj4ncI/f9/bzM6ddqCIAAbmJrTrwls4t39ec1DwhvrnPWhOORfW2mHCdAmX
mwdvXWwOHUM55rUJKdeOO112+prpK6XiT+jQHTqwvQLEquRffgATTpyS9n10B8TtYWuhjMn45bmi
QFaB3sFH6El8jZ2NL9LSrvZVP8FXoODvnI436vwKsrYrM9k7UHQ3IZk3yhsdxn0y0inDANhwyt7Z
VqqAQz3WvGDhH6liFZ8vcZRQ8m8eiSysgMNqi3lSMb5q1DsIXGHUJEbY9NKRbknys3yxJy+XgiNv
zW5FzOh3aOwETvHqaBwZXGbqPLXGmEDF8WAuMVIVJOpluiuyYTWVgbU0KqVzuqpaDIxXKTr6mTAK
hOAAP1Jt6Y/c+1Zq7sTgfFsGz5hS6zyOPx/2xR0srAg5GPYDF85ov+Gn4KvVBwy49LqdbuEMDIt9
eXwLv6aF2347fAr4dqZV5MMjHqB/smnOm8rTS+HGSVa9EL57Qibw85hnY1QZbBoJs6DRhdS0D/Ik
pEjArFZ33r/PMWnSjCbihzSw8bck3md1KqtVqaF2HYYV2DgyeK9P6CXSraPeRlPoV2Jo+P3MoyXG
NN0wsBK7w3YdAG5NnNdtksX08Drk2DvGNIZgBras8mtflfG2ko6dH2y27dEcvd3aUJHplR6osWib
1+oJAVLOBuWnOtNHilsNF2+4PV6akbyOHNFYo1jo4JA/ZntjSwb13HcbjItir9sJBFbeo4n7M7PO
WT/2YGNnoxpxSsKRuzkE3GXzY+rxRSVWo3Wu62zpYkA7kXE4VXa4Oc5Q/9NjNADunZEu9uy14148
3AvENnEyLzchjFwZRwet/7YQS+VIlbhikfGq3+jujF0F5eHXfvEp8zkugBVva0ZKaSOESPWpZ8Jb
o83cdnU+gkOpvvBEEGNYbb4bblZ2i1WX18BjqIa3Ygo/IVOwmX5+5elONJypLWhexDu6XWJn1JUQ
77sJAKLLOvXvSdVW8Q+fsr7FeH9Lr4ziOzm+ax23EVHjVLQxCIx7aHO8XqRngSKd2ZrTcQtowHT4
FORbgbeNTfhq2QHVVNX1M+omEVy0FN9FX1szjbbHriAYZnfBko9DF7G/LohGGMdof+ZhcPo/qvJm
QtikCZQGoJV6tBfuR4YldWbR9iy6Qlvv+sUf6DicKBi4kONaR2EaXw6hPmFZOvxeWfoWDzkorypt
sAQ823OqvoSi+CEhETjxdEevzXcj9Zx8fJfDnK8WBUqKV7JCE3SdPDJZCouC9dpCNSlnir+ZNvxV
dol8UTemwXkCAmdD8IkLQO68U0/kyV7Qp7ZUZeblDOR/U1Vsh7bxkLEXfimYHyvUqOfbdUU6Lpd6
/1+O0s7zpsXfJh6wYaRs5GTN2UICHLID8Js6POx1YGXroT6R4Am/ge9VUk9EkIOIy11bvmrZqTVu
Qyy1r4py4kxWa2fARPRvpwhjPaA7EfTlzf1DS5dSzN+aYQo9uL43RVGtrKjRZRlMDwSYPL005FiP
uoXO1nrZuPhmpLy2QbIIGEdZi3YvcC2dlq5g/GAYsEiccxL9mWn95WnT/LKsIKsGfcm8wQEzJLzy
V0bfGz3HGOmMxbFo4buR8Xm3msMw08pANVOHMSfIdy44t96ihwNkhvGAjVNhd8hvv01MsLEPbTZQ
zDOnNJnBA3srI9y4ZZdL1Q09jCZ7bLR5hH4EfEQR3DMKjIwrNjBLOIiKW1bfCFlxHPwJV8aEAhqQ
rJIuEKMXvFlS7Bje82AfJNpd/cU0THrE1ECbw8iWmBhVaJ5kiBWV7KZsjLTCmA2GzYj0/mHIF/RH
Zak39yep1kfmpNh3CBEtN42J+5x+BbKrUnL1CCjGmhGdG8Ai071jOyfWtUgpOSmNwmBWnP88vkrS
hg05n5MHJUh4q3EFkroAOUDlJ+fVbVsw4dT8ntOzvK3F9fPZ53Zbg/Pv4HsrHE/tFjUvrqDjfHi1
lu3eRaYdOJxas/4aMwrINbdyrZqs6oxVh6md93n8EoBQu9Ossvw4cD8xwsK5e1ID55JCYThX/idF
NjBV80dUCFVq3HlTnigil2qvatGo+cZKeF+C/aU7TSO/RvoYjWX2xjBZ/5RYl1eaupNhqadT5tZT
nhgb6EVFW6S5yewlv8SXgWWgjTPAfW/mB5C5grU1t3XJks8wGmjnGv3sJJnYj5NMCl1ujGygs/Ak
OHm1uAPx1HIm1/W34Duk9QMl+4iX3D3gnCRvzGh5fuxd6rnEwj8xmFLxcfrnZVQjiBz7VgQcxCQA
sDYqxKKN0dcXOgizqac4ooiJM7iboUWT9v5jV928lA+3hB+mwKP7K+ZYrThITgrsgZRo7BWwOm1r
zvVADG3yNdp4AwXRE8NeAow64war8gjwtH+TmPbMtHgEe2m9EA3Kq3OgNmmL+arADCvgIy4vxeiy
DLnqK1RqSSNDQ7oQuKVIwswy2ZCNm3YU2qiDBibfbTAUSjxHhTGlaGIy74Yrz4ALbWMlk854JZFa
34fRN9oyPMFiy8tc5McZYer11xjWcigB9X7k9T8dWx+yAIFMlAA+B9ilNGsuFhy8deNjsaXq3aFZ
/kfBt0lMT3Q9vr9rIzIMomVZmEbdHFUYgMt78DhfBoAVPGp2/jY1IiStMVKp2jJhLGt00Kvv2+n2
0KBai/AiIzWhu32Pl+xyjZuNTXUYQED3pGsHz0ILKHqF8poNWGlvRshE8mOLZwIeZXZInM7hsOPp
1hz14EGLe/9/jyLYcztJBSa6pKSrFTGMfx+r35QozdJWJjs/a3ABLV7o3JrMhS39Ni6pqEaGHPB9
M1CC26McdoL41lzSubUObcvaixtJe9knFH+F3RzAznnxEHI/V7CCjBwDzE3V3E9uHe4+zRqZHA6J
+lgEtCTaUoKcQK2rmTIGErByd4QoEJQIZLhSIMrDHnpC/8RMAu0i9w/l6461nvPZf5BVBu81GIxT
DcIDHvFhKS3X7C6fxG6SsdBmoYQmYYRIoPnsALVO6LCJTrC2wvTpP7oS5LSflvrCOXiKWyZPBM4M
u340rVTjDmxJO+4qjob4HPWgW0CiO//fufW7ewMl6y8ONXc1v4mOVTMvarLXBJ1Z7NlD/eFMcWha
nynenwSAjKsiB8LYIS8GYlQAAjSHbbupGtpoytFQjdJerCdfu93Na2jGW+RnsiIEgZ9MJCgIPNt3
DmkKrAmsUUz7v5VYfR1LYJdBS/nKFYr+YWGvQJdKo5Lu+aP3cvCOopKUfQMeExbPnFOaFy182kaX
hWDlyayJ1No5TKVKH8rVhypWgCnXL/ZysTMassPFdJB052e3ubndS0NGJU9L6T7oWuKF5opsLP5O
i91qw/8KqNHhELA/B1WBg3eAFhL+EFl0ocdRXDk+P2iOdJ+0mcmO60XxTzba0kx9u1RHJFitiUHZ
HWkDnHItAjCSo5s8qi6cq6HPJuNEncwoS2FNC/wMvlVxRueHhHO3BqfiygWADpMZvMBDmHkBYbEq
tYovnw6FJc+vEgXIzaI+lgsqPwza9IoYRmKYG0EGwIOtig+SX20s2M+gCO8DwehmpYrNqrMiIgpO
FFx4eN3rg+ataQ8ICRh9Y0p+e9K/L0KrIzb5Mkv9g7UHzovw7qC8o5c8s2Dkt/3oV2HJpQXMnVUL
xuJRVYR9MmndsbzvrmR3KyYimEtJONN14VmM1igBQj2FOtZ5aHYYUdDDFK9fk6l8NzOxkHhWlW05
jwAz0aEuSIqQFeEonYVRijhHUyLF8cHeT7yf99jR6B0JYgVHU7GCX7dVlhVQT/5ifSXH7hqbZA5T
G0swfu/29CTGBF37HjZaMeTaE/cM9KsCBUtk+nYdhsctc3b81EX7ZHqvkQN8xLd0mKZkBow2WYHn
Ir5HimNTYVK7nspSK6w7x0Mjr7G8D71o5TsHVQwI5HpVqPLnVHcD+Zgfs0kJs/b1o7K5vOYzMRaT
uMIePML4o4WXuJH1lf3QGYDpoFWcQkV9RfxDL9Wo/8eI8kWSq/Ry2pDjLoaqGunnMGkOW0Vht539
69DA5ksqGW0ooJAQe/hivI+XolpQbs7KhSu7DPISppOsDep9KEnJ7AUbASgql0535gi31hTOE2nH
7KHJPyEuLMNDB4h5jaZ+7XtmeYCHpYMgM4mXzcEjjVeRerFvOhXn9v8VwKCzChjFoVO3BkgnOl6B
iZCQCZv528RYJ0nPVsqEJLR5R3jGcg13mjfSNK3GdFdVNvw/SA1tXefaReoH00ekaRNlXwB5+GRZ
81+B7KCcmJo42g3ThofW78pjCQox8u9l68nkiuwRASj9hZmjnR8yGgsWuhDjdLR62OjlCKUPjs46
HvO0W/8oHEaECoxeHAsCB3wowwlT1ezTK1p+lxuo8AdUBrl7xioplTHsJRMqP68ydbRRkqV7RCtk
tDU2FpYCGU2Itkijt3FZTOCCJfAysZ3s2y2grq5mj8sywuK5kafo6JBKppZXj8Zdwalc9reej0vK
EQVax1bZFp+Aw+yNeetPfsC9I/tMUoPC3rcbIfJfaiBb8y/OaOPLSVBLsN9MTx/okJGWtxUlRFgR
a3FbWQ1u9sSMxM6+fw6uMIU++aR085htQRy1fc7NQJiyRaxzoL5qXmqxnTtlc/73WuKT64ZUpF2Q
Mqb1Hh3FIGytrWVkbyXNtfUdJdIgzC7j6c80wvaytzvl+xpoNpCMwlonD+T1cZIKcyI16rDNYJcR
2OjaUhcbkFYXmPa6ti1znXajj58PREjUsrfdwhCaICBvpYdfNp5Zr9cDVTXhlvF3BBKSHR9l/pep
8/kkkE+SneJLhO0kkfJY/IQxdA+yfLIgSOdt/ZyMdYBgB3636wJNUIVLpLkVSR0fKWhkZ2DCR3bB
Va8e+unPCzOmSb2/jcXgOOPEBEz1mjSr3BJ4ktcdV3pO6JhzFuztvvGVS7SAsADr3wTdW/wZU1I0
p95ciE3bQVWk4TQNOl7RbqoDt42PyTfJokncT/cUInprrF15VVxhddn0wvMfLahqA6ocu22z9c4D
XKZNuwvfBpbSntSePfiKP38gcBVHu3IwdjGwJM4ubjSGNrRJ6bnhB4c2eYzm9cNzTI4FptpIDaQ0
mK4p61E9aYwi/V06jdixEV+8XrcaF4SsDAlB7S16Ha++XE5/fuSzvRMIc2D5pdTKaw6tiJw1KSbG
Erl3BPACzmODQ+FbwCdq7ZTGsyd/L+K1gCdkqg6SsBAY6+Gcqsjhy+5YvK7W6ORUydnYmsYBn6Aw
LOg+cyIE4qPgFhU7ih3UHIlIL6XDuaPNoZRZzOuLjK3f8soeXuFNukEK8VthggI5BBfXvsW/ARDQ
/5l1s07ZDrtZB+W83E1tg/jDalI8LUOSw7n5KsjO4pwONT9xLe3e7Gx0pNvy2ZEbWmYZEFM62GY8
D0UllStEiXHmLXlddG8AbJ8YbL/3nzGtUh1iCPMgZUWty25RxF0AtM19IrEIaAVfV++bf4fSgO0M
cuf/HbzDja56+bE4Y6CpaS7FqKoCtT1vmOIv3HkA/5sGXQ4Cu0ZYEsQe4QOC1TNwO6LMgsY3AcQv
oz2XvB/MwFSt0F7tbPTeSkDGuQvzFPvAGfueuJxdCh4bVsEKnEqt1Sd+Sa/CbM3bBo/e63uXpPQA
7afjnzBNoNTsfPJrKb+UElpV9Q/g+eFNegpNxL+09OSrsBNVUp8zl1sh9ZZLUx7YUOJQfdZ6wQx3
n3U5U0mk7CwI1zxLX2UcMrN4mtAsYtUoR80t4s4GCE31YkmvkVx9zwmInNkUREyJgPWEZ+vXN3BZ
8LMpQU8Oqw8e7ek9kUWCyHnMJmOK2O/Elmjk5usR70TrOAA5zyCx9B3PasmIJxDZQ06HMF03dP2q
NtnNaB9051sPHpSQTCegRXKV+Lqy6Q/rkMAKCgKcQccf0ERcaxOypVpY1yycIYCMGSvf3RgcxbpY
wtfgRipU0LcY2Ly7KRcV5hjd7BurwsO2wnVdNjpFVHWxuiF5Bkdc/RlcX72XBu5MyFJqFk6b6T3P
9ZnbyA+3PkbQCnuvsGp5EJaBvDlbOX6BEkGPAKyBP+XwQ1VWKYX23qgocDdg1T9JHwSruUbX8pha
gZN82VeBCIej1bOXysItTmUme8EbhQdiuiN6IVqYfNVD1j2B7xWFvlgqdCHRwplRwJDYUDAc+hQ9
AP5GwXwpSrZIe/swur+o9Va84fjEHNAC0MZTtBU0ZPo+LK5ftO2v3i3/cXkZ3FLNq9/mMJW/NGmy
QZHhph/2i6S8MYOnThwg57cQ5zP4/mz0DMx/XyP6M59P3aeqUpWM4/TyZlo5L35oN2ITakPTqCfx
r3ff0WlXBX+QizjM1huBj4mp2R5Nutj4Q7aCee1zyhOYGayI38UNQm+dFent+Qjii8vNcHQy35Dz
cufFZMEx1St7kbWAMfzdht1T6T7M7MqiX6BV62C2MjD92F5ILhnTv6NGs/+exFOZY/yHP8gDATq8
kjqOcf9KJUdJTdnI1GxgsCToefo3r7YqkHUJ+NToN/GoG62a5RZ/hsEwkGX/jeeozCDV3LyuYP+F
JHmXvjkEFiCmfS8AZMr5KhJOCAH44LouBAp92Wxj2/URgkdpeogR+mina7J/C5DB4+Z7nBpJyqD2
RxWbEL1kSOSfY6PiPZ5eEIgBEva6Ub3meLtkN8uwJg6Sj/OU6CT9zq08rg7FfRYLbc1Os5A5jf9d
UeZxcrZ1jsQe9fKSfRl8/5wNnXu0hHKsRLkX0efaNXq5rePAVy7afCMAHbd6EE3jDZztsr2ZVGTj
q2ZcOLu51SKLd3lBSPB7HFcchr/EB8oooYHpk12Q9kFjUWN4pyMiF9tUByBRBtZ+JhbHORXE97ij
6C+wsYNugsI634DucVMfZolDoRxQodQlE2B23x94TIB9uNRKc2bwKOo1n9eBK9eLWmxD3u+gqSSx
sIe0SpYIPHPyqY9eDqePD1dEYccsB7a7/AeRo1vuGARegkSzNmii/DJ87NnIaBDMf3nHkD21TIhj
h8H7/tPZ3WzDZ7HzjQp/cbDc4xrsXkOz3hBNKS6uP1OcJR18BieWQ4hzkxav/if0Q3YBOn4ZogoY
lI1Sz3olrUt4QouhhbsrFYg3iLRss6Crls+uGYjXM3MTu/PQdJKM8x8LToA8/mfupQHLbsW6+p+E
9U1lZUKnVEaBX2cw7C33R7a9BNvJbuK66PuMKlaCUWs8v32HiLQx8A0SB8+Fw4Luk57SgV0hTrjn
Hu/eOLL0Bgu7slxmyyVHJ1hOXfpCN7k3B5k2YaACyyIbSIsBQhnI4+9lfkhHISmnGt0DdBblENKA
fAwl8A5bTjnsLhORyKmCNiupRTAZROmIhDaUD9pHzsVBeu9vW+X2oOsW0Ee/UCuoNPmlzrfdujjr
X1f2xunb0jDMmbtFfANP6esGuvqIAXW2MSmFMecE7zPV+fEShWLiy2S6daPBLuvowWX6w9fsfAr5
R5W6xowbyD637TC3zMkz0SgpJqTcgeCIpMWpBCG00LBsuMVn+pf6vWPBL8MvmOGb2hn1P9tp1PqW
eKmXLRcDqnBfJLwGYl2/0QCZ9KSCOfSYJSDZ6WmOcA8dfD+pasoTqpdMUOxDo5fRi/Wj06SYLkIz
UMljkO9l84U3/2g8jjUR3IlpjxmyT3uE6akPZ6FvXaFlx/gVAKj4jMeJF7U2U1a8cig06v1a/lJj
KSfpn1KP4OWUJtXvwZUyMYiJ6zNZnA1FUZntMu7YfvBU83onpQfQLOMNZ0cFTSPlOXUQb2QWwLfK
i2FOSdoldz1MZzTnxzqPO9u+R+9O0G4bRquE52cpojyyBxEy03N2+NwXsw9Q9uHYadwqMdrfPAqn
c5eQ76WgspKWZJVCSgAkxpfzdgyemOVkGv39UHGtn1mzUQ4TpctIu/Y2Wi8oS6NDoBkjsdBPvVV8
jpdMv7/jqMK0+mXzYj2Y6oipRNJM7cDCTDcF205PgETraJBRPuxh5r78B4e+I9C869xwTpqPAseD
zwHV9LvuHkHCRrgRBDuNHNJO+PX5NLIBDZVmWUOKlzPcZjbEa/Cvg0VnxsE/PxNmwx+QKAXQBjma
8Er6Xp0Vj+FUJ/hjHaTbQkCJHVT8lA9Md6oxiiIYgBXcJexby5ZgW7LjBOEi42T1TfO3cb/GtcxP
amcWSFf2ezHSPglEMCpDSCKkZ2VhKlhibsMbviHptEM0+bwUCUyxMQKHNs+UfFjay+7aSzj5FeiI
XW3IfxmSfQ3yLAFhB4L8DAhSUu5h032doJ9tXwU2FGUqUW5yqiJrQdX+uqvxwDtP4CSWntFqx69v
3WnaQGD0+VvDr/pY0LmCZalqq0FiJTPqlCKNp6wrarNyetG+6J2pLWWYTVTssovHUr6E/HcXWCTA
fQzn8PMWLfieUwojFT4zTPU9kxHR0BsYhw5F+bRDw7eKddgkVDzPYzX6PAFNYnmOZHlyixw7nsAQ
TZX3xV13ZyfFnFJbrkvyqQjSLshAZJC2wE9SUga1tfeJgBfuH9pq+pq1/zYmisy4p2YeYBiy+H3y
9afzSReR2Jm2PLIkz556BESDEwE7tHAR/nOioG2r4phbJhnYEBR0TcniimdJLLMl4CMAJyvpBWVA
wHjOktC+PRQZ0g8rXJfBoQwTp+aTYjtbNyy/e/Y69LzjaJ6GpSFW721cl9nHEsezIHy7Is0Y0mHG
rIfXOFyZfXEVnPK8WozuFWDLcYQEiXYaw28ogpTWOx5o3lpRAi2sYp5cKUPSMa0fowpeU/BPl4ch
lVdICI+eFWOkiAvM8747cv7lBp6yEdW5WqIaaludzlUnqGIDNkNbBJIxS3knG7TNHQTHe50p9slj
IJ1YNJ/nZoy+2cZYJ6tqV1GLw58G/D1cJO4/GEhhPu5ipJVLJWSIWMq5HNrPG1j5aZionvh7Y+Pm
q5Ugu4iy92LOniqP0tXfH3fgd2ZJ6+8vqACd2JUvDJWdSWNavvfcPVjPIopSotjiT5bFfpeAGJ5A
YEkDJFOeWCX7y7L9uyimWa2ReJgnvW7IlfAjtJdpj6efvNgX+GZbjuQwjNwXLIIzmZP8MhD0ulnJ
omh4c8O2wimQ/PlF6oTHAK+hfa4mcmEsfgYYlloUhAoIMOdouESXtBibx4n18/Lwn+Oco4QxVMhu
IATWM2Plt0nfe4z1fM8ltciDNwS8F1/+3zH1o7YYaaW+tFITZ+W2szYwGT0PMzDr6+b0ysUIUIpG
T7xU5P/EKkPwuIK4MLmUB4gq1hmw35PsKk0C/saME7F/4/FbuHnWc6TO1mNuAKktnl46Qd0XW7Ju
jifkRBgPme7RvBMfYYeDucffPNO7dQMbIhU6YLTxrTeFbB6tmMQPzoVGBF5WimBg3bktaoKU+O/S
xj1kHejV4HGiTWq2IzdtphBPqFhTzP48oDfEZ55Y/95DUxWDvyXsSjRZl6g6zg5AlXE3f+5/i2o9
VpMwT/hfzqoHOYLZ/cKlxGiUFl9gvy/cZ3bfKChWeM3EjpPbeManRtoVjM9JTy8DELL0/gldK7rN
pFkqjciximIjbZmiMeoCrND1QEM5+M/iZfuDw+DtB6V0B18+JbDJueSdYSr/CmCeYa/bdB3G074x
DGHD/YUlNDNX3WbMOaeLQI4P3dfpI5sH12KRCEo5bCM8kFsNzI9h/v+/29smOzUeXN43IgC+4JS2
a3d9VRlCwHO9C1eTM8FjV+sKrKKPvLwp062ef3ci7wt3x9bjjWlO6bvI9IbQZi8I+uVMNGVOTcGj
jIpqn1jnaY4FRGciQiSh+DWo1D7Hhspho6dZWCLzsvKrfqk5g//HrFkNAD7z/GN3asFe5L6u28kQ
Lyw5aT9CqrxnIwYrNZvSVJUTtleiqtAUoS7NtUBqhGvmio9uEYra9IyJrfYjMdm/WsjRJ97dB6U2
AEptZVLKwj6xn5A0yMtb9HY+eq7yXsK6S5RtGWn6vH5xGuUg56XUXlvqkpy7ODVc0Vx0yfwzBvxV
y9BSFKZWh10mh1aQ0Mm4E1HGo2FD6XgUegE2GpP3q25SU+EwWesdqCk2C0Glamqoxw3QJNsHDmoQ
t+2uMEto2Fkav4R29BK/UROK4nBP2onHFaGIS+/8U78b5pKwUopdjXFjeXqpLF6scF+8gszi+Ppr
jo0xK0DLRdRk+bU2HM/5G0z4DqKq6QoLjQXUxWjbkL+898eMhkVAe8+fYjsy8/bgcEN/JDffPEIx
5cZR/aUpCZH8pabPWFKBwtbaj2+ArUf8KSK61QhJzczCjTTlxeaykKuKlUfRGED52LDbrn2/3JC2
j/VQoagXUvG2CegUZ9wJOZmoLGpWbe7AzS5CQxFY6CPbqZgMuaw63AZU6RYe5rX0FoFTSARkylZM
yQZTjyVlMKcXVIhqw3XUPQstVL7ItYN1Wz6nK+1v1w+Vcq76JoEi7OE3fToKU0Vma3h5gfLu2HFm
mOzCzp5xvSV5qhad507g3TOLOvclwrc3hQfdjtystPyUzBo7mfBgEQdfIhjPrK0QrjLn6xaQfzsy
IRoLKFq8QkYqMjJ6X1FVr+oNF9Uyx5BpLcT7fnKEEKi/xPYd9YjceHDiC/6apKZk9iIg16SXRNpx
hqPdelaJMRy5RhkBm9lbT60W7TcbmXP8GTJaDB4QDCDTxeuwnGYjQ8cCOXbUkIpI5n4zPUHYegsK
cfZSD5z2WOTOnffaATHoEqZ2tv4LxMeRa/QLkkSOqdqSsUws7lTJuFEjrw2juJJIv04XtzYQof9b
Nmx5aWZZPMCAx8Vt2bVi3sULVl6ec1T8jiKVIA0DRhg8k7akS4iAEXvftTWedz/KXQZVHpHGNVyx
1OUiDfSsm/pxhi7AZDAX0QizBzFXQL/wIR3ESva1CBPL0mGdgE7XQUNYrvY1WuuMYCmrPvVFrt0a
rEKWmXsq5IaWqo/k+WNWX4O7re14X0MiWvbQNL8Ibk+ecDaM2opdS0HfrM2K/2K9cVXTWEDUmAJ9
A8UI5IRfTDaX5xqUOxHSTRYlHw84VBjAutzN3u3zlsBZilooq39bsVPdGCOiyoa1BAR5VkJfdk6m
D2QxrAI3ODjp6T0O4IH2EgwWEZPZXUW7fq9HoudRW5WFb9lg5+jvaAq04l6dQF5IuBk9tTfYEGTr
7OE/JiY6Y+7SGxDtkxfEy8Y+agJsc/lZ/3VmmAhrmdSD7cdZyc0wK2YQxEfy1ixHBtFNSlgaAekM
b+NJ5do2/V0BH4i4lRAgmA1+vTjcnYRBYRBT2s5h3UhiDOf4VofMtvaAmi2y/hzc+MUAdjFrj8ZW
JkR5JP++eSWtqzUJxUW2HxIW0hnd8aL/fhldcKAA4Y1wUNH7HwVa5Uc8GhGdCOHL7jQE3dvHwr1T
U83qyxFegoBfGLcO/IK3ZwLz7re9iTOHTKeFOhkEfyHUpKHB0UW/zOQA44JM6KoWYCpcOJC4FQ5U
XbftSpnh7xHSD4Qew9/AE6fjM99LusE4h7f7wLKXBer/+7kINICaGnrPDpBva4go325ZHJPRADd8
vIEmr12lg3OVbvExw+MDOeL0rCcgFa99Yz4PIXyl07BisosVDwvBzZEw/aO4f7eZPbI2wLSZpF5m
gVl4pkNdYogfWPfPS3n38t6vv5YXmE236Wi+T2p4tFaoafMTX1+GpHlGF6M8BKNeBxqF+8ABzH8B
ozZL70NNlg/R9hXMcXtEObt8VX+pYE7cWTgUWfK6/huIFdKRTY9/ls295fYCFBsZYES83yq8fASK
u43QsudQ3uDHm5oKnWFWWzEwDjlE8rhd3P8LbiYTEvg145WqqD5mSJF3TTZ8LdTXPqmODfCANFif
55RsUzgPN0bfchdEb4fmeQqxC9+zCAMXTIlucWImv+EDTzlT+Ld+j/baQUBFZkktMum4Z6jNDLZ5
FTkRc5Hf+cBVJZFupGH8l8rlanTHxhq8uzXS1ebKp8Z2ZyvnVUt96084j4f2nBF18DuMh+yQBNf1
QpQOyMBf2hXvg7JCmHpvyQ2LRvJWvHMAJHPndiPGdAXGbQeRgUPnOiwd7NDbgUIQr06+I08AHRU0
cefwXRNSq0jOXirgDNko4J9RSjT5gqXcTz9fPFQ0E0KgKFblugpfiTyXYjYqSBebW/9xAoJwBOw2
BR4YoD9lAvD3zwZiBwwGaY9K6k8zFJF6HWpYFDLgFISWG49gU8DkhzT35iyBdmgViPQZ5rqLbMv4
W9HTmpM1GUK0iMiRgrZYvx7iL2h3W0QiKZ8VyWf8tZ25eicYRRtZsdf/JiyZ1igfDIlTKoqSAB1P
PVUCIIRt7nXkLxSiFu8mJ4pXEl6wRi6Zq6zdUZNRCuMD2YccJiELeKjbw4cltS/vwDr62ayVtXvU
04aiOy8nb+CNSirKk5iDx5tj9Vn55b80DBbf+ts1CPrZknNnG3CS7/pNicBSSLDrGGoz3BCF0+Bz
3RR5dNnVBHlF63/haxH8INUTquFIyj5gryB8Z/JyQEa07k2VnUp4uoIw+u6SK/qBF/iORqYzZjHl
v4+ChCs1LS2pE7s7slqcbpYs6PXTgKL9p1h+FGr23fdLS7yDUGIEWAvR3yfRBD110kbyCIEgl5FQ
QImaY4hVAZ7VoILTULYgaJ9FWKAFXchC935xlU1V059pRmInABtU/QeCIaSwPKtmLJTE4GGQMSHY
/IEO73EDgmbh3wwWNiGmcN2AEFsKEO3/xvvsgY8nPjYxFDymG8XpUojJx6aP9fj6Z5pxnVZF6Srq
T8z4xE24agAyRRbXQ3+TT+/0angDaRn+xUApEwrGiwLD3giI6hcpYDrghy+ILEabTF3jPdbg/eYX
9N8j7WkMcO5+HmOWoLdU1/xSJzbv/oItZ3zeTyF+UgIANTaKM+r0aGdfBDa836XG1WHOZFULDgL6
KYexIhzCMlhDVqHzLk4x6WT/G/H/s2Ho68b+2DiGpuLbP8zdobQergtyIjnY4jivvtjdvJh/WowV
PfWX8NejWcUROqEaVUit9/LVPmUE7Q2yiCB5KodvCKC8gw71KYaBWS4KbPoDcxgZCYvx3CAXMxEe
LYV7gMdxAS5oK8MWhttne2mHZ8UV2RnBrnyZ5xt6FjKsjAVk0thTe4YbCe73O7Jn/yBleLYbcz2I
bHgUHcz3j8Q1Q4pe/5xGR9YCSOpdSV96WGpxkOgLWDTRlmXsizJQroGTiarPvbYKlqzG7QQo/qec
NCaZ2sVrhkYnZn6r75tbEN6uDj5w0MTygGDHLFxiFMrDrxGAhQiFtWMEtDOFVdMMqZUh3ivTgPgG
SYJMG8Q/5t0AlnVLhM1tDz6kAlqXn8LOkiSp65Cjx20t3bAW4VSZBGFr/l1hRNcBskOJ3rJR7WmO
G6idCiKO/C1DGvTHbrhEnmCxMndqY//TnGvNnoujpiBb96odgWCx/ACUR54X5G7NbTr+38vOOxhZ
TCGRqtkL3ljdLe0w4yb8eM34N/ZqzQv3rb8bzKxRWkbiSLgt/As+hn4HbmirtPdF/3u4i+kD5NLS
PDdMaCwO4ZdwuciJt7BfXBGbmiwkw7Kf9rD5NQEviPjO/DDUIZUUPkO4uiKHzWTd2BxSfE6/fyBi
h7jQ8hp01DQ97LM/bvLXpTs+GIrEY0FFSmXJRxElxnKvk9OL8ohnjw6Ku3oConSAM8s3xkcJ50dK
pngzj2qtSvEcSAKgLM64GPW4JuHVBOU0ESxehlIH/Hh25NKvLizwbKBamcU8Q+kNwE4xsvFGIdOE
8hqldT1vnxnec+kX+iHnTDlgeDXaldgknKmR+nBsp0FzDRKIdie6HUPhgVsrN6SRHvhpfeN8mgYX
XKQxnAKI8drOfxfQ4ck98aoXbmAfC/hf2ue+mxc4ZUVdww8ZF7pz/UyosuYeAvi24RUoJ0jGI7M8
gmefVtokwuKVxlGISjOTaGThQGyESEEYAicRor9V5ekS9iifndo3hNLFwxMfFCHFoNLzCLeEkAHs
/qjhj8mwAGy3ZqpsVAeI7KA+SAIweSn8dn9btcQg6QlHD+agUnPKW2Shz+PEitzsDjNhOnOvPyYS
Q6wbUTVuJhj+4zZ7WQ76xSp9H3i5JMv3zX0I4x3+nNC6bSPnKJOuV96cmdPSwo6yzsY53AfaUz4N
99uTgWjt4o2CfD9bhJJdCAO8nd+IwXCdPYG9eV5sgHqmkjtkkVLBpoZzk6ek/Xk8+M823UPEAwwo
XD2XiuRmXG8pkB/OS2Kmwk1DKmQgoKnZT8oXIwBY3aUc9rfmXshwPkiJnklcIpsIjEjRGpb71SIo
/BryxaPoOFMElXDR9R9RR3WguzMNO1GKBq2lbTulhHlAOfwPJ34Cr+I3+t1G7YLHwKPARTEFWS8X
xY3yyVAso4KGP5dpdw6INacpF+9pazIt1/B+dE9R8zgM+NgWHqKdieEhnrVoEdpvrdQlLh7kPQ7v
csFNeGXhaMoNt2tle8xup8vgORQURdunMXqHp50s3Rwv4tUs0aks9oDXqpaND3jmLAfM4iXsg405
hrZC+SugPWXUKbhCirEZ4XTvcw/FFYT24uQ3AqXT5jEsmXdjbjHKP3OnRj9MX9vYT1B/hetsY6kT
3tE47wzE3ZvoZTLr2LaqtYdkiMerYdmC/X5Hw4aJkew577O8+i7RaQZkaefaUn3SBdZdpbW+Gvnu
Du3IyTqbiyXf+IyYxHYIuA49HcuImmMAMnzY5cVRLVyIgzYb8d1l5UQGshqHuLSPriAdua8mYt2p
azcJpNHRUCiqbMHixmEiecg1xBqMsv4OU3rHErGiTFORhp9KI2OTFU3pzUTZuL8MVdKu23Quh1ki
GSxUx73qrTnF+gJkUMEKysMOadU8GwM+7W1LYEHkDHiVTbIVqe7jiLdsCnVyelqeMZgGDNjTwkT2
YCdeYqcKe006PwH71SQXL6Mt/rBIcyb2UxE0r8aDADX8T/Bsra+kfeAlRzgL4UNRd4oOIRbDCSun
RgRYs2S8j7076iv798GKBEToSTvIN6lH82bG+Ak9iURzaTf3cYhR7VDZAEvj+3omK/ZGhvaUnWQm
kY3Q8YHH7TLzLwdzc+AFMV5wAZ4OXqvtr+0pawKWR2d/JKsfmRJUS/3Dan/qWPnZH9iQdA3GwUa+
SDf3ewZb+pl/y4xaeh/R4e/F5N3q4UNgyuzSuPC3b28OnnHfW/RHsYTneHl/wxfBDFxgxSUhkh/V
v8j838K8maXFctEa6JiI/ltfCCxN+XDmt04yKzNlioCWVUV3YPha+rN9PwWd9wHKA0dH62sOO+bn
jMPYHb6V77avfPZKVWvpbEhQ6MEiQ7ConDGCKDlrcZMJhYal+WHfbRxK8Zmsg1O9Cq1pAKuRaQbp
cBslCi92ygLDzOwsfJZH7kQ0TaNQbb18eppieV4zTIzHE1Bif/3eYUEe2wX0EYI07neS/8RhwaTS
DaQxbnOaeR/5etJKVHgUKgIAmpz1dDncHSECRriOFBdzSq9lRcvZdsF516+8Ps9lQZ6CW8umqxyJ
XjjL2eGGMT48zpP3AZBg7mH2pm9HvHcAj1kmjZCtRr+DoBAJEVliwcZDyMF79G1LpL+W32SVfp6j
a5BLzxTfV1JKWXfRmu1CIVJo/u4r29wP7ctiypOQaXWufY/HyctrtShUmkrF/52Sn9LIM/dj2yVF
GwEsnIphITCkZ130OjZjVYoxBNounLbtg8sZzsk94eWV5maxlKxl2A2Ie6+Jedmq03Vryz9UClLt
PQ0ahpHPu9HasiSXOxe7Y5QPy3oL4UBOFoX1s3K5VE88h1WMarNgNXFsUoItBVSyDiZXJO2uMFSB
Hc0taRgLSLB2q7UuLZy1zhwFExacuiVds+zwIR6Kgs5IH2Ft2+mkY+CxuIpdOdMii0sy2RFLPXr8
LnovCgV5NrEDg1+sgRlovUIb+CPWrg7mS067PbOTFg+I86ecR5oh6Y8mBr0tSjLZlZMA9jOl0hp0
VXG6qdfftxN+zaNzOEaQodVVIdp57Fjz6o0rSB8Y4/6qgit9r3rH6BKiXn7WPxlPF+/9eZl+WXsy
t8LB+wKn+3ojbPtCK7ljGCHRbnhIVXfWcL8bhLhgyUjs45313JwdpK0xRhujtSpjtfORS4fsZFxf
+I+KfwzR1DTobnhqJ91WsdwlnfuMKMtMZgWmO0KWg0lOSCx7WtX28RqNr79cV0Zgh03mwEmKg5x7
Dg5G2E88I5Fsi+1dsH2MGA0Lg30BgHQ4M822jXV+ID5xQooEk1DasVDBbkrl4LjqOSmbcpM1dW5X
COgFSJicTkjIeZn/1OGwKCxDzCSzXadFPKqPsXg1f1da5hUwfIcuUBg6jf3qp5owu1OevWA2PVqM
sEK21NCGdXUco9ATehzgn5M4IB2kKSa+sX3PNHpe4WKNFfOcBv4ICCxy93cLCe83H7NjXLtrGOFi
LlPAhC73aHeUgRCf+bR6aWdxhf/zJi+GH+jFlfDNOvl36wOXgfBEaVkcxLHmQ4H1czbF18ZdJ6ri
WgRJ07ytfQ2wJxIL1N5e3YI6tccHjP62b70DS0mB5aYJ0j+jdhu/xRQTdk9Ok2qLgtfFKLZ5ixSP
zNqryJ4wZFRXmYvgmQxV8D3ciZHoRQYqW+T/VTyIIJx5a/MiK+opwsADn0e+jDw/1qtZK6QqiE49
0yWFcVZZBL+cupk6hsWXLknd+I+9HyQcmk/dYFh8Af9r4T0QMkijZ6E6fy353FdIhqiApZubzmwP
mVG7PVQbiC+MGH41qlX0wBYPC7VIPXwAKnnJAw1EKiI/hXQowe/CF9RXx+/5euDCE/EAREsaI6mr
tDU5I5Nze0Sj14eo/xa49iYcBytOkQZfAaiBQVLvNb+9+XNJvFmOJrF66i5NHjg2Z2R4lNG9nI9z
RMNLaoVJ/qh3OLhB3+zkCTAoAVEl+/73kLtZ8Pj9qIJZxI0N/VEwk7zKbeSGLrYBN6CsrfhATb2s
qV1csFCNOuWz7Yx7p46iqCyQJvjL6PC1e3GkYKy3NWpqf4fpvxI6nzncjZnoStzXuYtXrZu4SB2/
m4FzeZJP29pK94kRBAglGE1DBw+RYtcgMxB3Z1B3l+EYOz72ajmxjJgaIrrrSufu8E+S04MV68RH
1XJ/tV22lalC27ebHMgzV7jPfY0mjgaSssuGx0nwdGgtDenYjwvrrZAvZdVCuMsOK0dzMqYGzmuy
vmjFjCfLNQMukicImItJywwP7WFd2YhCgyESuhqIbT8YS9bAXoGgR0bXZ+zqw7IrsmrO+aCT6zG9
6LKRzRuUpJITOwquqmZmmL9RhejQhHmrQjLNBK81mVkl0iO4FiIcEORbedzxkurfJfqFvpesbIHh
gQsUaUyB/+0ZSKJ/pc59IuejRERCzYmpC25Tmg3r7544gXTg2qByr1JWXd+uy0RHtlVtQBkKJb6i
W2P4KQHlWXqldXsVgPavY1qHvgp423dbxGb001mqsw+H0Xku3GRuCcStlGLGx6wu270MtWc6694y
tfyj1b19aIs9eX8hFkHpMoN2xSJvKqzXnmfFJT38RKhmUpoSzupmX7Bmxgr3bU7okkL44SOxB3QI
lNnRr7hnIMoEuwPO60d10QYclSAh1p9YhEem1UIDRK/l8RronQbA5xQGOV8yj3JZgP6NjI55u2FX
Y8FzRs204E4SNf2z6cTyomI0l06MgMMQv7ci7iQmb7jsQEMqH1KhAq1gv/RXyYjn2chIWa2p7tZP
MC2wybyzLFLZSN12ezztcrFqLEA01VoOJWIHh+Flq3HJ7cqZsjzIjK962HYi1ZMQFVgRpoqmyfAi
5ylZOLBt3hPKs5je/qEtQRowAzF30N/T1iV0RAFkpb1j2kdBsmKObPJrAb6+mmxCAi6tuIsMdlH8
nDTaiEWCuSO6nYl7aw1TsdJ3xIBpqzqDHpKw7MRYapf1h4BaGVhqeHefPgN3BjnPRX82N+Cqtx7W
+Ja+JQJrch4tleQmEzxCKuM4oNAyBQ2ni1QQnAM1dji+gQ9AP93saBMWQwtQr0jJRHVklz/oUvkE
SDSra7NN3oPAKI/afvd9t/hnzsopxzXRrfuZXbTQYit4yh3GV5tDmIEJt7aPorQ7IOvGpRmgzvAQ
6W69lCMQbfSAoWJVk5RAPsYA027KJUuCDORH93UHyTTqDtcTU7W3X8j0Vsm4FzUWZXp2D/kZndLN
yIl0AeQjjZVV7/snh0be+Y/oOysEkeG8fctfigJpKT7P0PrdnjlZXHOFeDyosEV6DcHKp7+dBmII
kjv8McSUXf8VSdmyAf4SBvol3NIzWV5l6qWgHUuC6aLfdw1zHvwJXGYuQv1u7IHgF/f31q8bK5pk
ccvQYFmndf2jfoyNrA8oCHt/fz/+fxPro1X15cbS468deOpQcAAg7Gzhc1TQMocHxY4ZoBEFTBOy
QeGAELT+psa7numab0BkzPc1LEEcEGY3ldNGzlSyggfHU4i63XzQGsAmZvywB8JrpAATVN4TNeg7
4cgPrSq+B9A/VcD71ITo5UP/rSrhlb980z4/o3uUcHIUxXqPcG/Y7SveZTfIm8biJQBm0OusqJ2L
IsWXUH8Jjwz/+ofQFp5ghjASxeghjVDMMqxTtoLGaX+GPIGHkLwCEYTz1xOc8tP5RGk9oCnwFXdK
mzLjU0uI9tpVmS3yIyMehgV2Ij3FmsAGcPDzJynZUeJZZsMd0LTAPdIUDky/6yreJUp4zMUNeLy/
BSmEaFc7CGVeUcawooOqsxX60LXZ/oqvcpcH+BzceNaMjNWop6qH1MW8aIrF90NgnQ/QMAmpBGsR
A1ygqsy/Vps4zJ7SucXxAo3XeV0ze0Gvlov6jf6WXcjH6uqidvrbTPTaFmoIvAoT2lX7Bg0tDGOc
8vIi0kBK0+VurQf9AF3KLaqpFMGLa6scACrg1IrXNgRgIhe/otAZ+7PCeVye9GO/cc9PdWCVswQf
K00bMX9evR4YwU5qEDSuzQXQMUVI+xp+4f2AykFl6nmfw+IiUYOUUE7Rcmp5t7nxQVwYP1yKYPxo
BU3e98IdvouuFUREj0GcpTTfHE5MU4Aeo+sm5SMSTaWJUXZ0lth7L9MK7y6+sAc6r06g7Urnj3Sx
l6et3AKIYVYGhxbEdgKeeu5P4KOxSMybb9Pb3n2QZXtOw14iF0U7/84ngomlzsbEqgqTRikGXKdg
3gAUQF4bQdksPHIyUF1NZxJXHh3/R1HVQWB3qp8HyDzlWj3qeln74o3kjXvydknhmxqjhVm+GHEV
bXbl4kfAJ6ZuLJk7oi/6e9ejS21w0gTlc2FLU7uMdjdUrT9OtI8FvHDc+nt857B1Kj1g1Ogl3hrn
VBAPQIqUNF6l4nttz8wSqGe86yRvQmUZ6CsH/6Ifo+O3ciAaTLnWjqLhkmVlVdsHcLadG3ahizow
vszNfV62SEfyGQyheBPCrf6s1J1wO3HuqWYduo45tCoPzQzJAy9d3WVZREB39ptpsKm0Lc6PqmOm
c//Fl/XMjEYz0185HY30hkGD8HvdhDiYib+FxXraN+5Tw3cNITMacUYLGPjzIxha8XYbnfDnWF/P
XB5iAC6GxFNzkpcYE+4/hKp/9EeFUJXtHiPatgubCeoUgEQvpfKTWTVJXXTGR3gvEC3QYmZr0R8/
hB17EcGrc0wC3O+55eLjw9/9wMZ/kCZvA+RZ2pl9xBOz4xLWJGG7T8skhs+999u32ZBN+q9lGQBw
uE+TUKkpCBmVV2Oga+LkW4rRrQinmMmE35Ao2nARI/+5iYYqDwBz8SyUSxSLq9mnHkJ4sjOadvP+
od2SFxvAH/EjTURcsU6zrEm/d5O4/v+SlCUEBMqNHg0BEbeiHVYy5tSfl1oBhkTQzA3BRgWVxi4r
cz8Xp/pbidIWdicnJNzzrCuNGoy1nhfTj4tTQvJcPHGwvwS2ISIuV8IdzBSzqekTE6DBWPU5xCrR
+cEal908ti15KaHvoFOy5+gKRQa2UIjBh+Vnqea8VdT9kAC2ejvT3fbVSgr+pUC2ktMiUZKdAjaj
AMp0TQxfguD4my0oOaqFsk6Nl3dYQd0HytoSG71JeZuI211aXABsO2uBqzHAt4BFZ/oUk8r37vgi
QwoW2jHvxZ3UsReYEPy6FBctmwPerBl3OHcGqCxM3rMaf/nyD6datvhxk4kOCZQYClFZl7+FgSi3
KbC/m3usCMbg6+bZTHoW/YRhl1N6JNDdw/Psr1QhQffT5aSMzXAt1xDyhwyqD7qZrUPqvVDJBmJz
xhfmIegADA+untDq71TmK1Yn7CqYdy05yfobwQhxfCpO+WjpH03wJnG0/FrdzbwXjDpYgLxynVC6
YgBCAIyB4Tif1ZpcwULeRuEYplxevP9ingQwT7jrYvLeH2WvaERi5krk4K4HRWxq6nz9lrDCyw/V
4RK1RmEBYkfaXsIjjGCEG9+vFOr89UgzM4VkMgDUdQiCoUMLR+EprmZhVQ6FZD3w8QyQtDEyXrpU
kNReXE2ht6quF6GabWrGE0PuzVlEszpFuQ0z9zDHq31Lga6R5O9K7GpPhkET4SUW7Jz3A1SH1qZH
qPIShmqflCVSBUC2crYhXg7lKqhS8kExl2VtgxX1HWK7fBu5DmFXC1R6RB3GdlRFsQtlycXjTRD9
lq6gc21jp1FB85V7oUZZS2X1V9yT6cyRs5ML8QirlF7LzKHhs5M84YXeY4tgi4V5WRrGFwieqVhn
4Tpab0hH5JiP0mB27sa1ptegZm1pIgk/ZKRDsj5kbnEWHNBzgGkZXmKix4Cd0SaoAjrD3PbZJYXX
KPm/fSFz1RTCWDVzj5944m1/cFFKEfctcG6zUBue6qYt/tIMR4ZUtWcu7YSUfElM5GOPSOFrOzmS
J4wWYwSPYbMyLOmfHMFjm7WRKqXcgdeG52++E3wlRonR7VEejP4kqxr4oVLpyVoxfkVT1KdO10C9
6RBOt1jWvdSSGCe0ESBZPrz8Z/z/Ln4fImBP/jrPjE/kGu9l1ciNZfV5IJ03F7WyW1hkwLuOin+w
3X7TjUOgqi5ZYAJaq1PPZZ62arJ8dHFFlPtJNY9mZp3tIRjOh7JsKBcOp/EI8WE7JQCl0HUi96Qo
fqjkMBYzc541W2Gxe4GgkcNlR5CKH2K1q88dDp2FaRU5SXDYNyh83+X5XxUGecw8+y2b3Rzr0zoF
WjZBfMQVPglnUpUGjneBgQWTHmiX4aOuG3n0elU6ODYyBm4YescYRKfb22YqV89xxbJ11cPd9UmE
2wXsybvunC26nHnT2jeadTscnuGtcJvC8wWVA3uuUnAM4g+7uemua9xbmwB10OytV6vg5ONBA3hp
HU+bSTPf0ErTopFMrzRm8ztvL1Vs0ZlEHTKwJjfMgdZHxxcBTcpjSSR2k7nKOiRaRUu2McU6wsPg
N/2ibRU3tab6sgWge4aiBOoN9qoN3xdLeUOH9GUi9AC/CCWeBaanAWXrmbhvEQiDaPDGOjo4SQzR
ClpDQ1iY2ygSwTTGd0OuGXZeaeThS2R1SD7rdyEmwJXzLaWbv/0qig9cZ1NvSocN3QRF6scYaQFB
Sa7RS1XOXUf4n49UoaljtSlqcDBpYVgD0tUuj9qIFn6W7Mk89gVlxspg2E/5pAylIcBWxcZeXI4A
3v2cpMYIQRDiX7ekq44P6uM7oK/PYwbPpPVhH33M+5hGToxGYECzi5Xivx8OTiwZWmIAfmwy7Ba/
K8FvKzrOhYzLUYeK31JU8OC+unRI9NhlCSd/Ypw21D9NruKm2jnukRKNfY5bLDitNWMyScT0R6MF
VDieB1P0fCtdb+iLDnC4Cox+gxh258JlSslcs59oO/yqx5WIgK5zRhs7Yy0yooSqI464BV20rTcU
ft8r9d/3XTGT5zTq2nINmhFxWoShyiJ2fRY0bfFoxPgvryZQBIgSbzK0uXjB9U/RNyE18gfjDv3S
cVVTYJBEW1z8wei4EtlfoFP74zdiCaY8Ycg2+ZPjMhUZVJAGTuOtEzftjAR1KtzOoZMAFRt0jnpD
W6yfLtrCjKHFqI98B3nT8LyLD5WBoYmNMzI4BMcxdbdVpvIB8f5TiNEoPcDCGd3e5X/tFNVgs7Pv
mqBozv4NNhBNPu1iYbFsxLcN5vDMHBgZClE+PZVFX4xTBebbOooGbgSiJggOhXAisrkX0V+rmGdG
cT2lI+FSX0VRGgHwG8+7DKZlen+8MyELVecFd9YYubfvvFkylDRtTlDCbaTnlqc+8za6iU50BhWy
AMIhq9NjS1+Xofcwukio3eBHVTdd65DYTg7IU0+RDy4ZW01uDZRR09e8D/rnHNppGMCAccvyoi6a
5PzOwfQezZjvKMgS0H0c1ZNEyhbGzpTOPjSi9TlgzcY7mlrBxkhpzGiaqYhe5Huuc0W5ewUlSEZR
8bEjSDxmNr194p7IPGFUGKaGFo/fkbgqbmAm3rhIjatwQ1CjqmbmcMfycwW4Kn+hoo72OjLU0+YI
XBVJsKqmIquhSn2PV21P6hEhsYA3bKnRlyYLCv2yECngBt8dBUXHInF8UZJyaA4L7Swc3g2VXzAQ
Foxoz0xHqAMCBPiAdHYICJ/7InD7rk2n6nHe0gAWGQz9wc18MB46Fh4tbBqwbZSUuo/NaFo4Z3nZ
uZm4wVGKme3CT+Si3pncSbTpL1xymK35SWW8pE6/sLQDCAMBqlneX/OeupT23edL+KcfUbDnbkgC
UEsgz/bAi8gewpS6QzWYaPlDN1Xhwl0BZmJD9vgi2WnHF2hQOXz4xYnwcv6eDFAZjHdJQsNujGLV
plZjj8rvApvW5872i0c6aOLVujRbx4xitXct997szo7FR2HaGwVW50T+wyf0BVUbgk2yqqdOvN7u
KYVqFBGGLClNUcyMVD38FDEo5VM93SjksKTAHSL/3YkrsjmEoheyctjLybTcb/cHxgOUP7YqwNNo
/ef9tw+vzR16jPNv+iM0D6uS/NlSR2K/Q6G96mWGdN6wX51VqIGflf0fA6321Ev1QfhSVgxkW+z8
8Kt3mh1DkMzDX/8KDi+O3QBshBPxL57WA5cIu4IxObqa+AvFHF5wDHCR+0FGtU1uVxwau2pZOIUJ
lh9R0mMr5cPzbnwhttxhol6NeaC/R2vn5pH0gzOuIBv9eZR4kJamETz3Y4rBxZ+D9PyU8NElr5Az
IycMkjQMo744jfVvriMgz0S83gnS/M2KY4m6fKtcSIJ5EAXFP1FhXaegf3WFljKkKUgCHIZxanMV
X/TPUd5cfjkD7y9RPrLepRlU1tMGvGlrQcBJ2WJ0dZbCERhsTfPVaGhM+FicTA31jsWRTG3YK/dh
Yw3Q/l3ERgNVdpr/q4AX+xaFL2RJ/4BiLef9ZRNsxCeKvbpjOTjMEMkJe9vgpeBc1RxQTXj3udd/
4ukoPeUs1XnEyQ+vK44g3q2wyj9wztJmm27Iw+F7WfXWielbJuuRtSvlCzqEJ/zvMgEES/bVq1XT
lTOMGjKo7yJs/ctNXsS0wECVIF4JekkPrldFbKM6qsG5wFmzrW62AeOsCM1oBuhTV/WJYNB615sb
RKVIAQRUra5YurBiKVeVZIxs+rx7ZI1vdH+Ci61CkXMRbnh77nDbBHTsdf4pQS3Z7/4bqUrwqMbT
ZuAaDPH0GJFxgJpMRCedDlms4MhxHkkx38TDyjrdx2k2rWMtoj14Re1Jm6Qyr5yZvAj0qXX8xyyo
tsCH1dVQZ9TJDCI8VAYv9/clTI5Um7hGViqj03tmrbgq7M3gNJXgVbOIUgiJOaW87YmAUEreA5Ld
CGVuqY97mYFKAEh9HR0VDYWpH8h+mmCSM64IYHwo6hzu/SOCxJgLmzV2eA7HiJO9MYDnwNfrq1dz
ANsNM0+gb4FODIcfnfXN6VgkoEWx1Eh/obyjCqW24rTg6Fr/0odFe15kpMIETByuE5nOgy0UpV9t
mjkYik/9za/E2Dpv33qJaPtAmF5KMvs+uZoMmVg2mfLOpfl1IHcPgk/ZsU08lPeNwWcGu+v/C1RZ
57Z5XLxljS+s/ojmwascxLssJKp5oCeWBbECb8rY+I/EF7Mo2V9emErDHPcPhmnYpNyo20KwH79+
pS6en/FNWXwrhVuocgm1XXyw16lRvL1ZXjZ4p/w5eafir9KQ6ZrcQzYgSbi7vqpKUV1wd0WEOYcv
gt10+O47Ur7McFX1xAPR+JyfM9g3IXBXR0MbcfjYRNuz9DPNfa3qPshos5PQsHatG64acYpUhZXu
i9oRc4kcyqKpKkPxzT2e3kxZF99+LH1YxFBrVxQtCf15X+Iboj02jjx64xQewmiW3bilWMDU4fOu
YzrB3A9f+Oq4U1A9/BM/eqYHgd2q0KgNCmjYUTasNkG9N2CNLJkXmXdotMQnLlMSQWxnD0zvDMf3
6MV/CkUDGzwrPunlT3OFaff98SD9zVn9TMM5ummkky25C3eS9YRWJg8Durnd8Op92eWJF/CfW3f2
ozt7SFz1PRdjtm/wo80oRU1KmhLVlfMo0Iz7T6917LtBxtPiog3Tuk0s1CDdfXTlGtsxolzcQ3QO
LcjDj17y3zhvf/ZRDxUoU+CdNyBoLRTj6Cpg98w+MWsK3Ipzov0QZSTunxzf52jZqC8Df23X2QA+
CHl3BjXNNQ5frNfZNOdefgJw8NvH81/EyIWVH+t5NqnzSARzA+dAh1m5KM13aQ2miZKywGq+3vem
aE5FTs05Gy4O/8FumH4UkNqa61b3eXy/Ljr22byeQnh7J92FseGsqag+lAxcj/wOSP57nRJrViOU
x3wC1ScFyXcOoj7qhQPcKTyCU3FLmQMZtNX/66NhUAbhmfenUHLbWkFmAgUyYxoBSaJeOdVX3e7A
xYui4csGWEUvj2fRLx92lE5/xCCDAjw8oSdLvQ/VOBSD6AVZlJGfX0IxWHPFK1usk9pI/GR8KvnJ
Q/4oxCDvwjgSht/6xX4RtbX3lnKP8lDm+4GOmgJVfUsx0emHHa1FZq8NoHrht8t4iqmAY0xoN09Q
3+YLemjgmWtHv5NgGR6yLJsxKEpOh5L7dWLv/4ISwrd5maVmO14MJnpKTOOn7qMMCWrFMUdkt0jD
FSVvfPNh7DHMHcAb+QWjCxd2O3hVTUdew5Xi7Np8qYFLZRPvnaIaSAE8tXdH2JrsmMA75atWi1CC
7ZcJG+9dZh02YcA9M/CfEiNgJniludl/+X7Yav3q7doxrj7COdM5+C9EAhifXRi4QoOjZO/HZ8eu
vwlAPTQeybLHdLUzkq+bQaSBjqoNd5YLC32MzFVtNrVCemhsM99M2yPdhc7FaNZEynHhd9mFoMUx
l9sJUZpn547pN2+NA23CLtryfj4sVCDyxTovXlTSrxhRwhCaTOcfYM9W9Z+9GfVath5bjNNgzmBt
oF49/VnzkjhmqeB4hB/nFdXD+tQbXCZe6dHYodh5xi6hdlF5d2IWQ6bxfCyzY2S5OfEBoTHimhKj
FdWn5Iio2ixtFxPPNNtQ82EEMFMi0Eer2dhGa9sL3g1jh4dkiNUhudYS4XCZ1sio21qMJrjvsQ2O
d4dbPj1vFypwj2wwRbCLtm+oF7hoMN1TYjXzLV1pJxs9qnuGSnXN652IchBNiPEKCjXEyTLc19AP
dknITdifHJPGUCQ5lHtmAQTy+2aos9L9IUr0byyMvK0oRyIog3evv2hA01qMOsUNQFMIt1aAm2px
vppP84ZmOhRm5Rj15V+d9Bz7fgckox0CBK4wtTip6+L5HtGtyLFBwfA9sTS6qy5gDlHkWRN94GOJ
HM05Nh0WpGiGwP5ImHQ7gGu9CXBcr5V1yMl2+QX9sTz5Xw0mt7+VDMeN339a4RSR/53pw89Bzc8p
rXA/a1az7TikFuXeOA9IMIhYxUzyqrZAAsCplS29ordy30s68nS9DgPcKcZFvTMMAkI0zXsj5UaB
qEOSqxkzxUXeUycWh071JHw6BcRnhxkd1BDkC+actVJ/ikxa+oJsT4S5S4egG/BBzoUTEv3pP9ug
nRY+bxEyvmF2l6ZMxF5Q20NsAaq/9LFzN00gpK9ojjTEEtQmVJT/GfQBECFSERfwCtJ2jxmNXfBe
8TrU0uoOvLI+0viEuY7x/HdAisq11A8Nsby4LzutMs+ttQ76hkJ3q5AcQulcy8Znd1715N80C/Ei
8XEKJ3P/eKixPxMkfdZLtG2Kg2vKgqiKPzPtb5NDs4FBMNiwm1+ePiwj+Xc+fRmI7pSnhC3vvvMv
3RmupOVNtJ+Wv2G8k86el3MtnfNHSro/ylH0RXM4z0xvK1cr2gMDMOb7XJo8lkWlai9Potdg77k3
N9oeASHRuCdUYfUBRLLMiBVun+r+i8/1mjly1kahCZfj58XQ3zbFv8JVz2UGrCRzCDL9o46hyqaF
HPeyyARF++W8CSbwCFICsFBfai5ZDHhYOOe3Or4NKkIaqTROWgBmOmaGEVXmHywCVl+yPfRmVVeW
Hlfm2TMrivCs4tJOWQISupwZcquuqqcmlMDxIquRGX+LTs0Pq26QUCXGe/ngFkiteu60n9w5LNTS
Qk3HVl3/1YZ+jW1Z2gBXjGAqY/kwGG/Rb5jY0jSU1mmXdYGfw1I0Z+wWWVEK/ht3NaBEKK0PLOBK
aqxJEtcwntFNQf1gHG0Dl/w8k2ipxGTqsEuCYswvNi0S0uIyv3e5GvTf7kuDkYIqqJ01O0+nebZk
+UMgu4w7IHsIJYr2ydgZe+op8aECprY8NlWwzf+sGqml0z4vmpfwRPXtEC6oQs7DhSgx2ikStAMu
MxDr37ffSlbVGsUozN+/21tLLO8CuOIo7zJK/d3NgtPS1kAOXe9iF23Zv2PQ8+eS9WBKn2EW4HIO
3+C50yTUaO2Zq1JnqCo1k2GsJLtxPM40oDpm10JzjPozxAFF21W1EuGSOu4pI5uQ9MUBPvIsqlW1
ZSJsAl0/FAZfCVe8FwXwdwB5FN+zaO7f/yxKIxmkWy/pSC9RrNgcuUmv8UvDUD3TA8Q0u2MdUFzy
dzFI0i8Jn4j/8QENBVSueO6hvZCRLfjWiij2Tl3N5I/H/aMZaunXfswRGeCY2asTxfriMlIlDFm1
/EACIqedIglPkt43xtF4Kl33MvWP+CTLI//uyELoySXgKHDRoerKMzLkUMNqd4Dc7EOP9zZJ7x8F
GI8wJm054b6kj2VbwkkTMdv7rfKXVeVwXm0EKHqbdTYigxDmGpcIrCX7kFntyCcpt8Dp6jLctdpL
qkwLPWAxxZIe4YSc8Vk5N4HbYCd5h4uYNP4Jua+bE+MDtYs9aBjpK6eBFqf3Ksvnf8K4Qa+XY5/v
e7BbF1CpHW6VS5ATu7r7O7Qc+Pivp70aukA91J21ABKE6uhHumswjjpknRd4xF7pIcN7p9M/1OpL
/FfWLlfswDDrDoPu9yM5RnE6reytmO4QXhNyDabSYznMqre0SH9EwXjbNiA5K5fd6WdtXjbHNRdt
ib1M79dvikm8Z9JcK0RhuZmd3etmhXnWCeCeKL8I714XcgixRGZeEYdFn7L/mB5nuIljiieEaykF
TSpUQLsO9MwwHiFTO/+pjfeWvHrvRGv3DGAFAYeptTvMz0YCdLkCWodE46eDhI7b716KanC00+4K
NLz+ee21iEng5zYILLB5QzjEHIEQHnWt2knTGnjMS97JwF7clKtGDzapcDwoFQ4IUPhMeWXImSAY
babKiR9uLNF0oMJL771p+0F+lZw5VDubCKWzYR4bbn4Pc98bDCfg3Yi0nnMNcU4AbUg+zftvgSOt
UTc2OCiLIgeXFco+yyHVt2SXI/bR6W6FfRg1z6xV3lDbtpSI+jUTqBR5bE3WMQ3+csOnLhl3QzYM
N/L4bqiUztO/ErTynCooUUfU1MJBIcFsXi1zIPfujN6Ut5iVjKh/IwbvnjSO8NSdGghfl9VrZR2C
b6ElBi1jXLn8k9Bcpivja0Gsvh+oKEWel90u3IBkjFwF+YZGthReS4XcasquLl/s8/Q2eGHNIlES
PykcxBfDSFAXVZDLOGpBWa4R/1n8mh6bexZGNgUOb/ilBsp0MDhMs3q1yJ8zD6YHfbZyw2mDyBYO
8ydj3dXjcHdb7pqxWCh6SblCKtxUW5euLLE7fRNGNXbXG+5TQ5CqTVJqFJpB5dor/ZiBM/GvcIVr
FTBgWHJg9b7in60cj6Ysc3yF7WJbjhHFvCkP7WDjlprfAqCf0t8O87tdxRlf9bD7oSZtm3m+2i/6
SI+IwFy7CcfoIm5oF3T0BduFB6HgMODvvLQf5gCjHzgO6uM/wqfokQUNCHgEfusb6LVObQW63IDZ
V8msWjIwouHTPpI8jHRSzKDMbJK2mb7LntoUxAwn7/jrEn3rx8NcrMzvfy+LHZUmNAgdpDwPALEa
udTq9WnvT5b1WRzov6JVggfj1ucBg5SlxdJodKGOu42weQa29SVkOhPYbJyNzzzCURZ/RKol3Amb
Y3jpYaIWfc66kVPbAHeEWbKoq+DjihcWx7OZlYcIu5umIPH6iCnS812YNDczSpyniY2XbBjULcnW
rzVVUIazZN2n2Kc9aWhgVXHFTZid7oAry7FmjRMY76LFX8jiS1kIcbSzAcAq+O1jYIYORoF8sJIM
HSg63DMKbmd/o1dXgOscaHErqiUBYcK9xcvL8M2lSMQBR7GXXzc1YBW+oJ987Gy1WBXaAZxePjj+
tJXA5g0JSnlKkLYcEImvuzLznBI1lEBT6G//zHvs/fkOXms5OBcq9B4JvUr0JqJESFlE6ivrE/ek
ytBz6UqIUqztHkwOxDQvlMDzm1HG313VFvnRxEJUF9VY/s/279a9I1XUaNGqlHIRp4dRihxlf7ef
BVNFHRaGr1o5irJQHpebVVGa65tn4sN65hphAvDz8/E27fu4mRnI2KMFlt5VvpisYKy2fXWdZF3t
0n+hvO0vo5wis9pvx8USN5GggZuKuaos5CMuHimp7br6whRbb/twPz8cChzQYjoW+Yg1NSlMjRuW
2BlYs//ll7u/ifhi9R/pf0np+Kwf79wOFBdvNsIoA2vpHCtNWZDVfvcvfNEuixq5By1v++KdyCPj
qSK9iX4DgE0oZ6SOFrf8ihoITkU0nI1xlN11rQ4SLxO5ZPIqBvDHN7zWxEXgM6WhKqfDFmO0LYq0
7Mlcn+zBPdygXETCHSGDL0yJR/86nscyhAxluUdsboJmIcbuKk32YxOV0sVrQrK1SAuYhRwHz+DO
EM/MMXh0vr9vjQh8vBxAz7DGy8byyyspjmQJTB0Y1qxfh9NAUWRr7hx0yzo8d51je2k8k+5ABP7j
ilQpX7gocGaJekmSwEyuWcqB1YuuYW4J6mWHuiajDg7MI6GHhP1sHIgJswyUg1CEFD+Iu+07tDnz
WTzCh74Q/lG+xDJ3UHxqsQphugZ4Hqhzh0azkr9enO2qbHm6Li3klCNBk2hTled7CkQ57X62eFtx
vU/HoTbAqEjMkmRYdSXw85AvpV/9vn+czBtJpBLSwuexvYKv0EaOdNYn1PRDRU+BwcZqOBrLKD9D
hYvCOfpy8mU14k0HxlmkmmQiFPhxCH11dNYGuCixuSZW7q+YjgtKK2f/QdcbU+WvdwOhua6lvZG3
+rVxCi+OlbrfzCYI1s0JbvNzA3CfwagblU7CAsWJEP8EdA/01LncnTr2Vdw7VLE77k/pKMzWFJkh
5IxqB/PJl2yVZvfqpALJgp3rHGF0RwII9vRiWADcQQKoAkk8P7Me3RsKLwU9g09mZkMkiId2+uIg
VulDjK4qYfOgpvae2CdcLlgz4n8h6w5zfdw3qpOWU4XNl9EKWPvIPcop9e67JR1XyZ78qlLzCid7
NPhZlZsODKJXC2zUq+w0SBmAKbQdB5dCChlXrcEjoyMdHY7twQNnLref4NWWcwt9fXnQvbDaSpdw
PrLgrl0aA9y22emmoqZQteYOLv6KLzdPBT4El797w2AC9T2nY63iUC3nCyzAD/RshEZh8e50H44+
6QLru5PrjYN0Q7XN4giYKp5msNeq4i1zmET6zHSEyGI5hTdZ0kxQ19qMfNETdWEW0LfDh+y6mvCx
7nC+fr00hYYFWBZot9BjbuSRYoFF8jUR9g+Em7MdLaH+ah59/PZ/24JMIe5f5YAb8wSRIb81T3G5
6jn/1KtTgX1jiN2Z0B7LJ4qackzbiCPluo8GWFqifDO8igQRrB1YuKkpPxFRsAP3uCQrWBl0Hl9k
I26qptuYcHQwGRKCndecb+xoHpYbdTnWLvIkESysLrToZGkwKUnVJxQXx6yGRopA+rcCGXaBOJqP
FyKt4yimTChc5dfNy3lQoi3yhrz40ayvZyyPipGG/Oa4EyNmBZ8uq63YgJHybgfs0r3kKrfRmJF9
dtOdV2nyWXfvQUfBvnziRaTWt8NsKzjyMSTW/17BSOJ+osEcUaOs1KVt9HAQtfBXuonxPyRG4hdL
1lMVqECzkr/DFgHpw0Na+UJQd4saEWTOsVQLP21u4zFH87I4J0lQ1N6RIqX+IcdbCfICe8pDOqLc
XZK/jRYHMyCRG1VLM/TRSQyreGZox04MOX7bMoNcqQ4/rcEM8Ww7b4Qj+VUgsGnogtD7RvdN3EF8
lsW6NxajJsFs2ZapC4YkP3EDUvTFFSuZnkrm6XzndB7kUqDrA+sOZbusCWB+WdOb6C0F4JlJPZQc
SNjxGO2V/yfgItXvEE8SS4a0fVnbveFdjkK2QKZmxJjZsVlQHgzP+rt2gh95oD1BRl551FNQyqDl
NHfbwBl3hbZcDmFdnjDfzFuYeS33ubKUIt/jUx9WzsIjUDvWWY6CnJ4lGhc/FN1buG3IUk9ywQb0
MoeKrKeO84jXX18dosNn9onHBDMnC/BPwL8d5hP9xZL3YyKtvdgHxH6dq4XuC9NbfB9qQzSMXdk2
2exFbK2GOSzFhoWQDEeg63/B315Jwt/tljbqWk5LINApy1+7vwXu2MNkUaUvni2fKhKrKiJgR1xu
dzeHuJxAi2kSwFhbmWHR/AxDa5zWBsCcTDWnOuWbmyHHwj7cMAQ1uHKdrGntnm5bg6sJnbO+ksdk
4OfnFW6Lh4LMjGpETEC/GqEHx44N5XF7i2FpEvDoKnHULiDcB0FfXApNYOGAgpir1ENzy9VflYpM
t8Ai23YoGppGvapRvozMJQqisgnXKpo+8oefUyZAxlo/LzzpJxs4u6QWMgASu92vNIKjRgVlSnpS
b/HQig8s2aGexw3W98Md3DH2BXjbPHuC/OxsGw1f8SoAXr3MOTpphn2nEImYGWK8g+Xd7yuPFS+T
MYSq9snahVAk2KPvbUZGKp/agbOtLWY1ZvmYmbCLs6+xci6y4WFw14w+I3wrxsRJvTexCfycSv1C
KW7j/BYDR0ZpR7hBzwlpqsZcKbRRhU0EEQrZ2X5e2sOT/y8U2rLniL+NLYJBmFWx/hVGWpNF1bQY
6P4sEXlvNSKaeNH3C4Jtbjtazq1J4EFe6/+PIEyEQOLoNcFG8kpsFt3vk5kcjwNdNJk4ju5X/OnT
MohmSEQbmd4IEl5VdLeXUT0OQ2DY3VcIg1FHhNanfWYnwZuUvduKElmlo86lt6J+rwCxCWRIlydh
tUNm4Dzj6IjqVcwAZ6T1Dx1V6oy3wqoS4uJ6F8H/9AZ4eiSI/QBsDc+AcoFZSF2+HJnp6ZKKufRH
UmFD3IG6uvhXpAAbeLLCuhhXYQy5o5kkvAB81lS+VTcbnz7tIZi5yhVCZlJPOObAA9tAIUSMkh4M
sf6306DjQ6EiG9cyfgCRA1yLnUsMXTEXYZB1t80BxvzsxirL1XbirRirHXOxa+gWGnO5PvQ0dRwR
xnzMiCln0QXKYsHeQJlZwSMsYPCQTXbaUz3I7VQJD0SeOjgZSnTz4vyhr1/13e1TZCBWE6vBcFeY
cA7v2kNZz29TsjRfgSLJ+fIBTAL90Y4SqvTANcnZgyphAfwEZy2lxihzw0UYOHDuDVIDClUq36FE
PvigshGr4RE5JwZ/GufZ6FGl1qgmhu7jfLttVZ4eRCpkwgPOUctiJh+yca7oyY4x6CFRh79oC5AJ
t2rrsnzPHIriqNTeWhhRrQiBH7xG0bU15viKI1SANnZtHb6mRBMwgJrogkHIQuoiTuoyhs/oRXY8
BN87cgvCYXI8er1l2cAXszXFgQ4nrEDYpPgH9pUNHDiFK3gegxxt/fE7cuCU69zsXmhmTv9jC1Js
e8n7KhVQGkYQk7acYP40RkNS4vXlQJ/gLwVX2Om85bX0ro80kSs2fGZHWN+f41BD+wUnWwH3JG7i
bQd0LDy7I9pxsCflWXXL3oQeDtxcX5qD8Njm+fVasahGxK0oER1+YLtIjlxwPK4odygw7mQpJn9D
7s+IfZxLDD6+BzZpQbl3DAvUEJu6rgdcApBi0XGTwDJKR/I27kZySCJTAMejLdoj/ykkUARO+YmS
FQ+CwR6YpeWiDBBRfxT79pwPTS7soopuZD9hKh5lO7rDt+HFisM+BO9NrfVxmSS57fNsigSYPXGt
neZuncYoX99Vt5dCG2Tjwvaca2YYXiwAow1fDb7IdZLHcF8TdAQ/rMkXCUSGdG+eTd+D265HYwiq
2BaIMIpsgbR4CJ8KeTDUNx+RgEgZ+Q62SdgAiDUlpT49VovH2k173PSkSxLzlw/IQxYDyFHY9mtc
Dh9sDZbdPdoM7sosdXvJJqBt74qebKjCpknl9JDxY1oJ52RPfakf8ThJYWnmrmkYk6c+6kCrEWyb
BQLDJwCqwkQBhwpIPuLxPsXG+C+HTFWs7u2uXbapCo10OSeQX/zzenQB1n7UFxWsXNLRhsmbkYnb
ddkddNtv3kJ/emg4HeQgxOGgrL8ZLSX6sXVqJeuBD9vSA1iSeWF3KzHzyDcfzMWQdk0mlPqZBHvy
PE92ZKPL8NYsK1uhCUwm0+hztMqkIrjOSUhncgWwV0CKjnjeUzwRGfnmSKlSQVbKcOPJWYl9oLH9
vtB/v1rMtNUKprOCSKla+qZWNgWkfM9bfA6noxwbHcwPriQiteiMZ9p5wNF0KfeE08N3Zjj6lENU
j+ZXsYoQr+/DuQV8VldEZVdQ5gCIMFsrsTuQlKXxhs/p6OsQIJdxxIPnbukhm6Ky2cuXEygB6iGh
cW9IAsUPBQ2j1WKNURDJjYD9KJnlSjUF5pwOZW33smLYWkE9VIt8zGPsGjhl0nObnKcim2Lg285O
AvSQXj7DX3JmDKzyWM+xNYAS66yTFnlK76iG9V3u3K6IbbRm9WjnsNqyQzrlifV2W2ncIF2aYFBn
vkZy5S/Ji9ILzgv40vTfUyEFvY2kZ/hJBF8opGDDa1G/dnYZUh4x/OEPzeUJtFRRlXfW1uLuAxxJ
2PIodpJWEnoWatlfSqh7sPXPfMK7o6ha5aXL5KrKmLcQ24rTyNy90+qhq5VJ+//QP4XFd8mTwx5B
ElMfcPe1LEGYxF5dCTMnIOuD5WCbGAz8388l+MF6ZCMlnfhfh9B+l2GgSDrsAwEPJ9vtqldKiv8N
iKv8qdxZh0GzPzleaHLxqhR+11Vfm+Cm+6FWGHVDlPYr19gzbrkMrJD5cFZhcrXVQs1QhR5qVuyV
XZopulIbhX3jynWYJjLvR5cSSsEIjgz0LIpC13LNfzgE3WdjiFX8ubPkRLx3wuogB0ehCdB3su1f
SAkObLJ24DMDWauyk1drJ/Eq9VHmdANrP5xtwlZBkQ7q6hwAJBrYZQXdVnpX+rn+Ez06RsqatF4a
SzzjXdFSHyxH2bgZfDNup7/P9xbuCGioM6HppifmaKojHtdNUdsCNKh6ra6AKIZLYyTmPYCT1iwC
DBzkBNZmkOigU0zAa5Ay5IpjDphNrHVLeailxY+VXLcSIXryKOwGehYBDJ4QNhW8fuEwQIqZymRA
hwFZamzUwj2CuZ2MXXgD9AfdnG2FVzmgKwf1enGKUxCTzqS+5/XUhV5ODrkmL40goiaff33US5M6
aHBIqZzsgv7xGKIxA11HMQ+YV+S4K2kSPX2zmf4KuRLZan8+uT3VeRqOCFkKM0LWpxeKp3+xTRg+
mDbBmChlNX8EhtloiHALP396+zlyPvlaWuZNVkX4J7O5oCHJ1x5XO+Ib72c/59HHUYXaTdFBSmB5
Z+1fuN+llgYPM0q2K7MEJQSKqJfM0wG4S1Lbl88ykhv79kQdpl+Z/DhjWAalcGnJMVr6C74yKnVE
NFoZLTp1p8NgcH/+pAJvfKHKAzP3rX4QkuB4U2qu+fSvMJTgabilM21ktR6wDeFLHb1uD/b9mJ0R
dKysJhMT4ndCeJi3WqxfNN2SxFttQbT6bZZaSflCj2OaCb3tzXjm6Dkywjo9LGMW2Pu2iWsIFTIA
dO6z1xpoBWYj8ZNgLlSN8KLyb5J2s28ehpki600WFffP5r81AoxVIYxYBEtn7jK8zymnqfmM2yVB
h564Ux8E1MwM3NCAGGaj+IqrdA/cWfAvqyYbyQGuxt+Xp3kLX2aHhLTtmvVboe1UYmtDu8j9AvLB
2oS1zn1pM1gvGqW+r8uI8U34UHTPEDm0PJO0E3XaFbtVzmU7+rQsEAFIczx9Si084s5xJgs9wyHK
yykXJztMHce+wiC97NBzRtKDE25ZxYQrAXRY8W7gym4/I+81IW/Bqcg5AMWUuZ7nwMTbkfYXMdiC
RtZfCPF/fjF6obC4qznIPQz4o5V+egFjt16TCGg3VNfUHf1Kxft4RQAIzTrpEtmIZBw4lXms8GTd
B/0oo+uZgCvqKWOme15RYIqFwu0y00YK1VFFaMz0RD48BhA0oCfeUL56rtU/fpK3U95xLI5f5D7s
rTcmr6+Mcuwx0Cgzg4v1G+UUxOXvFbJ/niueUu++9YQivDvxNeseEzXn9N4DtA10Pl1Evjydn8hT
/KiukhXuHiISwtltrisasnRQDB4mBlz+C71GxUGyqJFQBuijskM+vzVxkgjhxGW8wVtenE2L5U2G
3P1u7T9MM1rn0CemCPH4wkwxH6lOjiMadMK4R4uxlmb5DEXWWn0q7WijKxdXahOvgVb+9T77VUe1
I8JQCQdq/VaiQR6qOFozUu+xxGvewm0Ui5SfKLojshplLYqH1bkyMIj8ayED4vhCiXxSfbRGpxIP
a1C3ny3oW8pFzBnxpl9EytNJwgt0Ax6QN2Tk+rr37LhJbwHnKmKRWCmQrAWc8JD/L4jewKj0rBid
Rb4ISGMJC1/M72LWPxYWmLlnRYo6ISb51/bWgRQhPcB575opN8VYrMFLWC6E0x1iSZ/qUx3Iymvt
BR+od8yyz2cKdCgbOBQDrkSGS6EP2n3yinmpo+kF2z/vVHMd8fOI7iLE7ST21nayKhnonA+a+OFn
ex7IckNj66yufxH6KPzMMq3zzmqrId2tlxq58zuJXzrMo+6bfLa6QNq11JlSe0YF8JciXgxo0G/s
Sv3xy1V+6i7C7LStcG+mSjVfVgTxVsZrip86K9W5uLblnwqLwjAOnDVor9A6kySX/QsOby29wLo6
eSRwQrPVQ9/KNavtO/mKHZWkLNqH/q86coOXq4uPRHZmOZ+Z6AMHhOqXj0qeWg6GnHsnvz4UnyvE
WKaAJsC03Xtw6L8qAeHHSTOPU3urWvYPHQqZolOMm5Rx8Qk6IFFUfNc+z/J9aPqVgOpQbWY94YKD
jlGaF4bKyPH6EciFqARFo+Z0/gEyY0Etwfq7+vHic5vkTfA0rCSC8HoY9RZ1/qK2PAn5d7LVMSJ1
FjbWJqrsnEt1+kAeTk3PFW/cNKNDJK+X3TH5iEHA0cqitLQQLxHqZ1m7wxBgMXRTiObz1y0+Y/xV
OFqL1k94nyLeptrjuwx4qg53RaIXSvkNQVKVUOBBPBEHoM0SHQKh7kZ1Cb99Iq/Pw01zFnloy+3p
3gVXNpDM1Lbomft79xPO3pKcEIuAA348+ZcVkQHAlYowPhl8qz6fBpjMotbE8a+N1lbT5iyb3a5U
VYYctXXi0SckSggENH/8AGKNR4cx5hEh28pFe5GVm44AsGBySdP70Vg5mqGzFfWM1dhpFGjpv+Jr
8j8ue4QFiIfKKyLb8scO60meWEBpi1AM+VCL0jEeit4EYtoiFydcm15SRuuWZ6J5ia44pHJ8ju2I
4V6uNaagIEKcQZL2+8ZfM13VClwYnIptkhld+q2krrlZosBJMroKSembXeewff79h0pUNqQh2mlY
4jb2nQYvu7D6NytLXoyzxx+TbRe3gagizkF3SBRV/oOmXwmIsEjyxKLKFkQEb7ZwfjT7gi1ZMnt8
KtQqvAGmuxIttxXxS7IXQWOrYOOc7qcTyvuZfNummMW8I5r0FbQufJ1fa1KEU+8uv76qfRbo6k5y
yqxhC4IpwqjJm9Wdzvj5HguuZBPeCXhbiWCcJHBe2jILw+NzTjqaLmSbdZemq+/KTm0W01oogFOo
2J1bf4x+gOQOQ68CvhjNAx70LSrO4+sNCwYJa6phvEQYci7lWPp96OBD0L1aBJJO+S8QomQ0KvnL
3ZoWVd3zPLqOVGxAoVr0ok+xsU47U3ruF3eFKJ/snfGmkU3WsStF5YnZLAvShqEMZEuXSKN0GU2R
lWSHWHY4+oHxmsko86dkmtwatbrynJvwKr9xGxLMvXVAq5OmH07TNr5oUzPuf3diXKralSMpelRX
sJL+fmUQobUkgsN5Z5p5JOfNWQb5dLlEyhgos3NUCi2MOu3m8/xr68yrqNekZpHsIVgJjhjQHQyh
EmjU+KuZLIt5SA6RaOEI2Y2HB16aa3LHP+gMeoh7v7v9MjIYur3A73uFV7l2CeJ5m90U231aFq+Z
fMTv/e5VahC44iNHfPVPssihOmojNL3UijnDZhMksi2k8DFkQ9JbeamgS4QuebCyuTPH+HGlheho
C9tvKbdYB5hDqMViSNWG8rbjWgcZSVICfdahfSm6wK9lDub11OKpxOKxlAO1XIbzveTo4UWIeyDJ
Ea8bZHFAO8Sd1l3Uz7N8aEKc0a/aa6HUEVrOGrpS/GzQukjEgd+W7AnpJCAAJEsRuQC2rU7Jm+DZ
WIX8eBBqUR8xD/EiLZOToBhUv2byubBCujHPp69D6ORkG0w+B5buAgLWjYyDp8iTXjF7L5sbDqvF
kdM1K+IuaRgrPOEoqVrq0jhrdQEWaMoO47OCKUMaM5DE9FnuB0mj76nTITAKJ4ZI89iffaVksqiN
QS1ljlAml61daxxeoeOEydbPBfeDmfYaGPTynA2Zv6EE+k3r/Sk2fpzazT04l8aRqOH1H0Z+z9kx
anMszgXdYidlu0hU58h320srBHVuvLEjEERRQBPo+DcujbCwCOFNVO09MN0EUmk8dh0hP5KmhGA+
wA+YO/3MHikFaLiy0df/vCyjNFKm3qFWN0G9FVqMrt+URH9lonyL/OznF2JkfXXp/yB8vHrN6AXa
KptWwyspMUkjHK9XDyW272wMwvJ0Sooq+crSCUYoaUom8+A1JyTDmrSupxfoGnXsLrYwGoKIk8vD
Wvc/RC6MNBgho9YbHXyZCgwm1Zx1qj17qkHV0xGZBhxEyjZHFiIo/mZBqGi27nHWsxDQqJr2m+oS
tTquIYynj9eP+oXt54ncHc2a36NUNyoL5IztdP9RucZLRqVeQJDtvCXmEoaMLbf1ZBpVFNaTRqEW
zd1UlOg8hUSaMW9CpqJlKpnQSdqUpI7UKWdte/qDG7mY6lr+/TRFtQ3Cr2ZGDUaPbxkLsjiaMxPY
M2kEC71i/jsDqEpCL5CAPWzMpanHxv4/mQWW3CArJ4KSivmY1oRmAVF0Ohej8Yu9jrPe0iMqmwr/
zWEFkLcX2QmDwCnZiUvQ6KpX65ECfnIM5nHlamKCvn13CDVuomfTq2vkVhFMwhHiqcxcqPCSrdlD
k7feZ2VaT3Evpit5otjrvYCAlZJFJ4NwIGkYO82u0cErTYiy5Om2jnASfEfsV0h3AjFAqq3zOypf
bepf4Ful9xv1vhyEzQ8QRmM5zBkcF0rYlDVpg+3abXJAGDQR4VMLL9ZWCkpIwYgXA222Lqmx56h5
sNwNXn2pOcKd6gc0hoztyWFmPGjSRwbR2K46pjdq7VRFFweYPmk4TvbQ86Ko9eowrqwTuam5CDbg
diW5Ek7H8dEyOIcnL+ODF3+j+nmx1MP3RoZ1ZlydLZl+6fMvDQT7QUjfSerTZ+fPUqpv6Wjbx601
jSMqGxZhdNLK5Xy5C09wqaCfxQXfIzxL+sEJkjUe/nwcnIXQ9aylnyirimxk+hvSNeDox9bmpKaS
PWsvBRiZ+4Lh6AwsvPEFMVF+wstwcwCA1IPRBGjhvHXXfuwXXWm1s8NvVGdEbm1AI4t/f4Sjfbkl
TicTlJKRUvMwEbu1wqpoavoHUH1lKkdGKQyOs43euAlNnZerlwsX33ZuvIPWlymtSP8G5xAfbiQ3
WC8ujVDdBWON+DES0xUk1p8p/wVFUy7ikTJSoIFg7h9VR8x72PmI3KSW0tzvVFdKAsHkSwAituvw
LLw0VqqQqJ5pvNw5/dqxILOpWfod1/XxW8YX2m8OU/tVqyBu8Dwrmtj/+xMNe2NVdZk996Rik2m0
2aBdpSVPDfkxERjueAov4xXN8hJC0F7L4c1Z9QiAzqZNY/0XT4DF99XnS5KGE/bV8Gd+Df+mGzKd
9tLNdd94Cwz+MfTsgcwoNuRHqCoha37llg1Qaq3w9NyR86BWTfqq6OO8+7818a8efjulj9bH+CTb
If41vSseNmaAaHjkFyxigsj094otTkNrmK3io7taQk2j0DeGfghip9QEHg43AUM2z1GlshgDArRS
tPNuC6UeFBrqwSmevJxfZ0ftqw1C81FF9xW2CgoUcyScUdHlhhZeFZDMKb2t16l4NEk10LNo+bRp
Drt5tiE1zwG8lshlzAXCHxjGqXkG8T8nYjgDslQOLzNd564DjOaxjTIsh6cbcs0RoKA1ZXQxNJcd
yT6tlZAoXwnZm+vV6dso+9GDWwPZJgvQj39PZy9KdwhYvO8T/UFrlieyRkN0ABS5gje37QKGYXrx
VMrp9Nsg60rdNDG5F/ijnHodrj2/QMZWILmR68ef1w+CJE4rFOcG3o00a6E3w/UOqJCV2GtsQhDz
wkcRLetJvs7oloWsyXlFBvx+czFG25+WzyDRwhlmubhenT9ig+CJpG7/yCcASSVYTJX7rN1xAQss
RyNSXyzB5HEMwQDc0cWEdljIP4F7vPygKSf2tmaQ9jdCbVDza/vgAZ5TB1sJ5ym2SJdzfGpjjUz0
yoq/icp+aYCXelmc1WrcKch8VQwCcMOoUNEM5P0SXIIGiJ1Fhcp5PH+OX4EQBl17lzDRe+hcA8JY
chalwrEUmMc7J2vIvY3OmSkjQFw5J+oYQVcwO5CKciS/HCSuawhyCMl0Taerac3ta6jQ74I4LBmG
4h1oXJbks/MC+FGegfFGoiszbo0drNul/zYQUwzsstc5O2sGauMPrskpT/r5XamyEHDlq8opSusY
V52W+tgHQDXnxyd+SactAZipXHgRvWapeP43hBk/2ZPmVocA8bo/wYHdb0kulDw/DMIbU1VMd4tW
aj9WObuwMZ7bNB/UkXWhI4CrfEnzU3+hL7sI8GYDUergXR2JsVDXw+RDmptYd66PM9nAFVf0G6Hn
QAM0uiWZs9F/XK/6Lfj/y55m4BAeYtfYZApI+ou/z9qS+XskuZkZxy01taRmxYTAZgDyfqFtquPK
+I2gbQlgin2sTvFDqddAq3b3r1JcCnaXmRCTd1iTd0WJCKY6NNiE4x5rswZ0G5M20oYlxQR1brgh
tnpD1OtpO3KkeCff2rUWHgJnp5Ym4z8Ey8bYNPzcz1wpqDkkSxSI06bYGaWgGXzpOFTsyvz7Vh9W
FfXygfn0BW0YB7hCNMbD3aMkJaulg/36C8OyUMv/mqhnLLW/2lp6//zALVWt8R7zakSIidkkkwqU
N+btk+2pBiP3T18ai0yb5qKMc3+TrIih9c68j5szqq2XWig8PBrnWFhGL09NNhowPpjkkUG69t28
h1/4czxIIJUjWgVvBi5iwsWsFRJfaZ7QkzzZRbxZUTw4NNfNJIi7i/GljJLBCjfGJndFG/CL521p
9uS7X6XJ1uyToupc9SWXn1+JLGfDRfVU/4+j3mfojfOlGfULSg5Hmfb2PO2Y4PomwqJrYgUAmLyv
/L/5Oy6FBCKoDu/6nRfw8wmpZqdk3hvZPC7yuVCAa0yLPpYsn7E/DIb/VWBaJRFBLgZydyMILmK4
I/bYLuYoEzoQrDoKM0A/3ub/U3zcRsvFGhpcEboswse5uDvAs2/8rK9kO8+h1POWL//AUn8QBBR1
UnqXpEh1b2Brj1uIgKXCBsXq9ws90mh6f01rXNPHfsZ086u8DBLK4gCu4W540OXNGes3UpRu1L+x
uXjPK6aVVXVpb8EOW3x+LW+2ER7MaaAWzoycDiol2doL+6w7Uci+Nig3/iLwVM3BNjTNP+4nmE/Z
o4BC0lCm+Gsy1eryUxnA2mHQ33cygnqgyAtYlFoYVyvccWSvxD5L0frgT/0uCV/SDxfWJtLkbkvO
3CsUrccX7hwwM+162EHn3+IiWRteluteFNkpFHAZv67er/YVTvQoVoe8HzTAhyKnfx4rdxifZcF6
EIJOASm4PI3W1avZJrZHIe6IbmHqdXsEj0ESuzzf+wxFt7ELKQ5p1tGRRQ/TiEQe+uzyrorMKjXe
/9dk8NAbgoW3I3aq5cDOQ8Q0znWxAW+ZNAMsHltJc9UOCJUsBDvtp5QAejPdYCJn4EqAciBbUpMh
RM8ShpsxVXew4ebZKtEZs6TKhSb/C7vMy7WGEibGI9rkMoN1l+5dYMsOJB3fy64vlhHc9w7t3mMk
9iF6/ceZaLiTbSky+wvviT1ZHX4mUPELKWApzu43Am7BpkaCneoizJpwm10iQGCykDhHG9JAVKJl
roA9q1VULD9iXmNEmeownvroTYdyJpo9pyzvqLn5dadrD93LsBUpufV66EdrH5Gq1R/TyrHlblhK
fh+vSebdNEWTsFZmnDtiaOOlLV8QcdKTbS4rBqj4Ef5O+pLwf/ZXu47kFu+RlJBgT4tzuTo7bHnL
GsJnPdXpaLonHCBQddia3D7s7FL/uVbp1KNCeVT0bjDWjYNfJjAPPaSnJ9w8yZsJa4y6qg6D40IK
XevI5/7D3A5xjyfFHAUpWazAM813bmiURniASZDPUBE1LaMV/Q7xMhPIhhIMJplpGjXXoLdY+GtY
Vnk2uPxCscLxxL4YQvXhbMryKw9Y0ou4iifqC8fC3PL9gNAjvpAFKCDuUsKMEhgYb8da9TLnsy6h
hSQ8/n1vYGGtoF+U6xbDr3or5uw9sH9LmzORBxHHp5JlWxyLVzDziw7t9hZTX7PW8mshk3Rpx59a
aetwLFI+eDh33VGkWVZRZa512aRKjaRX3S19aCrnsCjikuXRqguFE4p06EK67Ioc6IXN6LQM4DQ9
AhGxWONNKip8imgVveOp9VAX3QF2KTh0Dz8AQv9E9JoxmpERvh3xJL3miqEfuAJoOAj3dDWVhAik
0XL3R0O8vu/wFEctENgCBmPgFlZua4AvOhNzjLkLoDuU25YnYMF/P4IHA325BTSyJjrv9vafsJin
2N4rtUc0cRpCBqkenSCQhmQ1Qqap2Xk4pGkFAXh/+3MnbBj1CDoA4MYg1OD7oShLKTri+Pv206e0
Y5O/hBDihHGBnEfzoEnmo2YE/PirnEOFlA8zggsdDuhXEqLNvl9hhJSSniHc/ep10TidiLvNwyaI
mVIjmmwgru2b5werW/Dy+G0PAT+dlXUt8zT4DYJPAAMmdLBV+6hJEEhhfTOelH/WCINFPGfTPcC+
XaJuVzYaie8e27u+rUN3FnzyQPS9LvJP6ydXFaQjXdRefAbFr4OG48Yd5AyX8mVNfoYMCJ9XbBdU
k1SHOqE5BGay8LFV/QvlLzaX5ppTGXWFJacr7st/9MpGAOgov3IkA2QipFVh7tHlOGvV88y9eBlx
+Xuw2/ePkbKzx5tBNterzImDv9+BoKp2GiPVacx2s1klWYV8jamJo3e4hVg64HLJ+2TzlTQpwvOU
lvqyzozBPws7KyVcaPc/DjYK/CvQzMnkz486Tl45lkDq+JQv9X42GSu8pVTca+84kmzgaPH8+4Jw
qMX5fDgXxT12cGjlvgCduS4eFCTj7GRhlbpvCWNKdHz6ugnj8JsSWL71TOZQelWioO0Yji2mE7Jd
KgtB9Ay4QJQq1sXfj6ly6xYM1djr/i0oyyHFWoXcX5aXOwapR+Cex9GuZFTprReSj2eaioNzyuvv
vZazALGcIk7JnzSb4m3RXRuKYsBOiTe2Aao/IKF4K360mtnJZyeOaeFi6nt5nICZq3QWyx4BrVEM
33Vyn0LRsRH8xLrapfGuPmSiFnvHxd1QlqFTLKIx2jr2O0vAo3H+G8hpqvNu8hTevY/q2uiZEWaK
eRRdzQR3+6RKPeESGmEwmTYz9QFdPfsFs+RDY837PuFm1+TaKH0Q4pSEEuZ4m/k+emfek9PwNLWm
NqZrdKmjJ97gKIxTS04NFKHmhrHQcx1NSvBaye4gs3ED5EX5EdbwwkycTVoqxFB7ixCR+0T3RSOz
d9bNZVTMNtwtFRuwag39NCr88BmtizB4sw11AWRUaBL1g7U1O7yvLXv/oEpBmS2Ld7VDJQPLHF8L
15fjV2OS0s06WPoppkb8n/AJxSHlDjqU6fUUrUuhrKFjEFaN7R8u0Cbpew0AIsGfVUDUM0oG3j+f
BvTPxFY4b859CaiwOUjMLwYIHvKvEp3f33+eZNzr/d6bP9R05e1LieijcE9hBdjaA0VMF7Ldp51C
oBxp0sH6X3vDqloeDqdy+YsHRK2rtE2XIKFPkZHC6I1XFNH/4ahn7w95cX1ZSK3r1Kd6xQK84nNY
xlyU1bvPtaGMXzkarMwM6tj9y3T7buuNTkDbePNb18i8euBGOwEfmdCtfYNb2zeeXBm6fqm7da2B
kI1HpO1zkoRPdeg4wNg5mVlgum8ePRp1ocD8DH2div8ynnKbLC6cDEiLymcW59+9NG6jr1NLCtjr
M0/T2BEVzVqW0FOTE0h32cn6Oq70dLEJdz6pOfD093pYnq9DqVKH3nue2QkDpZdOQfLwXrUA/AgQ
W2Xlr8gApiLB5UlGGxgwLk9kVA3EnAwxZ03MXEXgJq1FH4u4C0YI4cQKlJGE7kHH77o0KZR99XuL
f66xaMV4E13nI59Axf0fCFeriHP9jqrrzNhQmwzuw2fXo3wa6nXW2g3Ft950rFi3jZfqZRDMvfTh
BUOV80rZGV6UWTgLoE+RHWnyGXiQKVWMb3T8Jjc8Aox5gOyZMzVmTT/2b6Epdb/6qzqVwJd5xVWq
HstV8mS+BjB6AgQp2rMSfOpPXAD7Yux+Zlu2XeF7uuao+hKmUJwhV0FsQZCbwPWsYNlK7BAfzG+K
ZAkUnQUwoTAeQbzVUpMw0uwMkRB/cQxidFlMY/V8OTfHeCbEzvVCTC8FMVzRuQjEQf6uruxXkMLb
OEuYFJH7NmCzDqxFj/gfjv1VWHwb/6ITUJdnxBsWp/eCkSxjw+akg9slEmxfzcMKu/VapUUIx5Cz
qKiuU521p1I461ZmSwsMUHddGteI2IA1Wli+/qulq0u4r2uh6k1Hb7b5u4AtVyxxFPz66dSuL6/a
WZM2soNAqbIioBg95/FSsDiDHqQEYmlr7D/E3x/rxf/WYZ5tgRq3F0griE5BV/3mOZcZ6yivI+jM
ppof3+FiyrE1PGSTqyR6x05MgYU8lnTScQI+ShpvDQ0t5kD2ad8Ft5VCu13dP4TVVOiqCtl/aPm8
lYpVOJng4e4hR9kbAyw51x/vo9lS4u/U41ZCTZTG+hHtseFPc1eUys3UcRntp5BnhqKHmn/tR08P
XyUKZcldOzJasX70nbciO2x8IBUD9hvQghbdj3qzP4tXiY8kKIHW9XyCWaj68KmQI05Dn3Uoa08w
tZwEXZsRsAzV37VWaCi8yyvzcvSyJTXRLfM8yY66G5c3Iog27bTmfAiTwga2Op7oTSL9gEpN7VmQ
3go7xrJCHViSV7qi1bs9Lc7zezubpsIoNveGWMqzeVKhSF3Leq2E+VsAHKAHBCQh/3osdfK4U8/F
Eiu5cdTDQYPs8W/5Pkhr5CcK1mQ+97VNv47/vYBHJwQFU3IR077Gs7bTLUI07ehQNGaxUSjvSR1Z
yUswWVUhjYUBFVDpi/vH1d/EBg/HN/2E1pGOLsn087ESfjw0qXl8DHnoyOulE8PfzLGp+Sr0AxcT
4wucIEUN89vNtEk0aX1fa3k+vceHg6v83qbWM3bPbDBTvxATGdDmOg7SSg4aHADxPnFIZC+4Kf/S
DoSgO7jnM1OCVTqOQZ+VctVuhN8lMZim7ueEN7+JSTDrhjsJtiaHkLEKfK/1z+tMygTnJq31pmbp
XLDJZa8b3LkHc+sOh6pVuS6cSLMyVYPbnVqsf8hokJjK67MouFUv+gf1RAFB/0AC+PO0TrCB1jpd
FyDM+v03zaQgKlPDAD5qC1o0vU7hwqeQdKGfTeD53azn6yMQNcmKsJyZ9T6rggGVb3bmQ0gfuVG+
2ZiGdqUb74VHDUihxjeLizhmBxvRtqBacdzhDSFrjZ393RNhB0Ruo2pNsWuVYXBDBmCdCsDO68d/
l8VQUNDMLgIdkSkyPvurtECaZ2X7hGZOohTZDjBDCFN/jY7TzWE2S0X0POcsWE2GUfVAqTYf9YzT
FfASrfSiewlYW8OjAxzcqyoSO9Le0aTXkL7c8JNd0H3rFqcvweik9443zhzHvYCoHViPqLo6WG88
VvlMJqe7/gc/IT/hE9bJb2liex1Q2g2aM4xHM1maYJI9SLR5ufoxneG3ABBNXOqWDn2Gl2/5e32H
tzsGSMx4/PGZArCn/Q6U3AvDbLch8D3XaNxs3lGSbteZkmoNppg7TAiYv0QyLAPttmlu6O//VX1l
CwX+TCvZ8YseG2/RKgAtCVVWkbuRM+gQXZk3Q4WXVsoBkfGW7LeG3PubSALepGNdiN8kaz7Y0PRo
6YgF+JTbu91/T2klkUiytBNUKKiIPXV3q3oHuONOdJj41KEOQiT6KKHqhVM5zrlRC7RQwC55xnG0
ewNzO9CG2/v8SwopgnT81w1wnI1Uu4W0aiBm5hv6Zp0Hh0P/FTm360xdjWPd/fhOhntmtuG+wiSy
3Hv3mdZbbcoEQBLkodeSD50s2hqefMbSWtXbq5w/EgiOdnSfBcSoreHQQYUb9iCFkIozIT+k9zd/
QzeELYp+j/oDa51gT2sO5ZgtbFEJ3yapO6o+UTh0Z0QW4GxjIMlIeMPbcdBfmDNDvuWvrabmzyjL
O/ODysP6YiPgztK07waXEAldIDox6oYgW307uhBblnV7EozzwuQO4fgurkrLfpyojaKrdsDlT+6N
m0/65zaLuj2gn8dPtc4Mhd4pQQI71TIsxAlI0PnfD7Pr7x6Cdpr53yR/XrM/XTOFElpFlXAvyejE
jB7PR0E2TPpAq4YlMZZBhlURYPPREKAUX9b2i57XaTrCZI2KxJnj0VhSCGRLH6FjweBn34JmUvlr
gY5eW5buTOCdyEIEPgecD0iYM/qYIZrV/5qV+gS6VAtWfET1hvYk30FNJcWGPF6ls6yr9ndL6keZ
/n7wid5WMomgNhWKKKl4BIvmsDR+vB+9gdSeXS2202bAXxi3t8yM5EEtkRKg9/Bt4w/d0ckTQiKl
3rmLOtamq57FNI0mOGadGm4V5lSmPZqQpgfEbRotHLtvlAw/fYQKhM1xiNYTzINSUXSwnlHVLJka
aDsXLYNfCJLKqaYqA40XjjmdkcEJdTbhdu8/TTlaY9nJ9zdV5c+56LCpoaoJXbvBmn0v7fUFtqUm
95kftXLdZTiHK/TgVJ7h64M7xDpxe+ybcGixtRuGFX4FfGHVkSHDOf36R27HQyCkQysvJj8EG+SA
+sqW1QmqhpTWoyRpFY41sTENHkfGX7fiTdfGqKfYX4C8o4rwFpj2P5O/XQb0CAhrcht5zOqTNg80
H6oPCZ3S1x5huhGd8b1pwvn4fOjz7WjfTGOqnmzb7AxQoUKfbD7hqSRqQfopCLDglSgIs/IeVkIo
YDNI5AIgPCFQHuySMxTwt3rhc7d3fNFX8IXsbh8k54dRnPg36ywWsajMi1dQl+7dWXFhCbN+grqc
W+DwcMcJiQFUerKtOeylt9HtSjefxbAEnHwE8s8NRjf4y1clWJHsVKDH2P9w1JPyA/YMFARga6+g
y6jtFJM4+DFvtDtu7MBuqbzcRYkDq+nhlbYaYevj1fFtcBxMsVORiH2hkRoUysjSQZ1EegaGueoP
6adNiD+tUpaGc/bl6NZ/Nb96oI9PhC+R5/0HaP5ceueU3xnZyVaoZw1ctm2tlzfhrjqCD5ZJq0ZN
SV5q6Nk2zstUVh3b4wGmM971l31ZLkreLsJdao+EZj70aUX0hW9nqEdW7DIPZonBoYZnSd2aHpME
BfjQZx7iQbOmYPoYvmh6LzRN/vgPXvhhsiHsd5EcVQJUGV5b16qDsrkMcd3M3NgHDMACifVguapg
hMgfYNxDHNTa8c76mtHFsb2lyJXweio4fook2GbDtXaM6aMf26BNj3Lnh+BATeKvZSYQRrlNIPJ9
BfUDIa5QTBiIg7qQYxT8zETjlBqaX+fkKLuoI7L8tJ2NQB7xV07rjRG0wgz5uyU/tT70VvMAzdnV
cyg9aQs+kNO7AfmLlA7rPf1O8ewjAMqrSEgUQhMdrwOHPhZcNOdr6jx36t1HkleIIVWuzFcesNTB
58Bo3lioMLEmgubQSNtARfFCJfiiHLKOB4YcXzFhAj2yHNaMI5lvHeC+tucXqk58T15250OpY0QN
fcmYqutfGjO0N5qgnbhCWh/gGaKb5n8bOVNUM2QSGaf2yRFhagKtBuOcJhu+BQFfsdyhVYY64r3A
ZsAYZaLMFDq7XkDdV6fRNV2DQmU5JoOFXJ7TGT5tXAMtcfhX6W7xAQLGcmVutngN5IZ4qLJ+5hxz
yVyrUvx2IFsDz031aLKVJXnAyi5WC4V7MBzvKFRt+N1LAaFVYKy4C21HCMcWyU1Zy8OvaeaU2SMO
zoiuDK8v8jz23VOQTXKR7jYDguiygG4AYc3/SzB2nUazPeerNryzpQPVCsyc8nxLDT9swYltY7wp
Jjbe1BtFJWLBVjZrz5b6Ffs8RRti5RuEYBGMrsCuF4cmgh5tmrzaWeIUrTj8HoeDqPYlEgflF6s3
JXhMsRiZnfAd8Ea4SblpY331Cq/2+jD7G/yrtmfmjMMbOKXZVGq7ESkz3vtTez+IIyXJv0y72v1k
C6hfriaRir9de7ADBXmFJBN58JyWuxR8wilnD4Zqwn2C+QDA6eW6OGV//jvTh5gSjtJuVMisL9PX
KDULp6kLWvwIwcJO0KVm5668ypoJZL/W43NGBMuKy/ROzPpzGXDxp3HNkTb24c5NlTRSJRd9Rht9
Q//B6MPFXAj4E7+U7PfFChAYTQ28Kg3Ce2NnNn+k1pFYAQtetawnytWWhDwVL3RLuagmunOUeZVs
EzSUMZhVs48vR6OIeDNbwSVPa/e5JvaDNKDXZo6acdy6lr+6Hh+tKWMz+y1GOMPERCxzykPF7kFT
9ost2a34mt0xMey4esXUvBCL6vJ8OEqNT5xssz39TQOZBzVqtMEjHmkfitF1esWeR6+IrRNOtzIo
aEtaFtU2m2SLifRkwEWmMdpimw6W3fq5PPALGdzOkGwTudP5876biQeLzFlOfzXW8SaZACcOpEHi
h9thipr4rsJl0gSARuWry10HsqbaDsETu8q/6qzHoBN1r5qxfliOG6SMmNmHTWtU7JMXvk7+Hyd8
s5exvk1hcUochO2xehI1i6mrZeiBy3lNAo7wO68Wfj2/HDSlLGKby2RTwXfC8mUf6z9CnHfUpNov
kKg5UJHSoL9YN3EpjtN/ekWbIPlA9on9J9irvh1mGQEGUjMUw7F5KVwZ+ClXFoOMDtk1T36ehPb0
ijGCpL7/py3VRxmOL1ZlCh0w33NaFGuejn5b5utxhRcV35BUhJ822Vl7EWr9BoVVkkC2GS1caZBE
AQObEc4rz/C73TALP/pDYRCorGcjcZfMHlthyzctPdIIM3hkYpX2BMxyG/6aesyHYeVyJag11dxH
BKEr79y9VXEsZ6fS7cR+PnYlX84+ylWgqSJFGwfOK+sWSHdEsGWpoPsRn+7KmqAWsycITvd/sBJA
80B9PBIgKU7/NaKAIECGLZ5jr0G29UK2o3Vbf0yqw2O9cNaxJ3awtJqGf8+gqgwVC1VH/VmfKIpc
EgJYJehFvz8ZjHsIilHy6iTqxjRY/GuWkiiC+XpNlq7LfIKYBFp9k6TYFr92EigaXsUluJb69BnQ
cMQS5vSMrwmNRT0fFmaQUWRiH015osEIN4EoNr5uf+kdAIHI1ua+YEg7CWepA2PlmgPIIF14Cq3i
MsJ79qVEYxsUb7O+u3n7DqbIwZPTWCf6FsdRaaokXgVe7yyx/cFgTEocDEwM6cokxI6seL3NwctW
kbEO7OJRoz3oSrLi07jsXNim3neZJy5ogEMAM4I7TASnT3SzwNoJ9ZSuHC433MQQjurFPe0ODBvS
yVbloKeOX8r5E1+T6HR8iSFXDvaxoPoHUg93aombIjQKP3cuVmxJI+WKpq0AscOh0xwKWdDth9gB
fY1hHmkejEO7hbn8R8FPrH3XnY3xrz0kR0hsc+wfmuh7iSZ46Hnnz1xIFVG0KMGNw0IB98aMUczO
gXxbiLSSH6xcFzgMQwXvLUQhh3HZMOayM1tDgVoXjuFaRGyDgzeoZGgu8DfpORWoDuqewG/LtjF7
+D2xWsUjHzcDG1+68qYQg0SIYjnEECmZcq/YToYAhu/K3Bh7wtRFIz2AcHZoo11sJzkK2gsRP9ZB
Nt6L9snXEYukUaNebMQd1ro6i2LQa3AIL8OAZVjob1dp5ewxJLbK01Lu4kCF+sNrFIj4SBM1xIhC
v718J05irVNtrUzlcfw2gRg6KEWN9GVI5rfDEsv2znQoi0rVmxRVEruz0Q6pewoYGPgtf5Q0dC0y
m4mCW0TQMWlhztffy3UcK9UjQynjP9SpcT/Wy45vurgeYOuDroxiAis1ZlK4PbP8G1ZDJqQfjFkR
+CRpE/sup3MegfoSVXcF6JML3lViNK/5NYFsnuchtRi/JckT0D6t7Ve11YcDdGrjWiu4U1lTrNX7
rDwa28ozQmyR0vsIkskjC8SgilUN9HtkWgyx8eoCKGeqiX4J/JI7B59XkNUhxiTt1mNDV0J6fxLm
5xoklDNQQt2OFouLZ+GRecpBi+yV68yljBqJBMHGdWZ3sccgb2NL6zQ9WLrQ0k72yMF85+SHGFd6
kpoWahdqoa7XbTNA/jQ7YicPRzDUU0ESP+V8jy3lSWQ9bHwSZgyrCnRrdX0SXq2MrNbUUASL0G0Y
RVhRc7iFNv752s7iW1dq0xPewD6uJHHvYb2MP3COxi8Lk/wvMzI3qcAY7NkpsjUcRnCoq7cU7scF
7s3CXoCDqUuPE2H6cy9W5s+9GWXUNLVy7zKr33h9qVmwSJJVscmV35BbtHTbHG9dnLhVZ3zI0rqW
bP7ywh7yA0lcFQiXUpdH0XWvI4O7U4L+Bd7gbAELvCaLIb5oj9rDGpRRxNfm7AlRFgmy/GDWjAog
w5DA+A1ysFXzV/6pBYNvpoD0jJIF98l8ut+CQZs+/5voOwg3NsngsFJgHpUfdvbhYdtTpE6qJZ5b
abRgDe/4Fe3YpAtKTNB9ZcEqA0bghxhraGGE68UxJrRdRUPXjFoQaXch/6OYVu/0FzNc7cgOlkhx
XKVEO1lawtXCz5GPzKi1F8585co1GDp0ZqFkCh1/nrJrhvOUu0aMFgzVBOlsFdiDzyV+EwKZUzQc
i8RpuUraWHDtPeCSucbFE+PjFlza2OtPYsWBuon1uScn4bJJdG4t4dZNkVvwxRVlbK2lQuXrPUIa
+ubRkLdbEij4HJpIhU752/kj4VOvpHwuhsqMDBtNA/aGczaUWLCq3G81eIjtXr68q084PsOSJ0JV
JbusI+HpP94uFLXI/cT6+rB4J3kQ20Ar32o8FC7Wzyutk/uCctOTKIdOMWw1FLHlemqiesOyKV+f
9az6mB5dnoEBJ6qqMyKLgNp4jgxz5av1s6igQ2Vii0XzueeLyV52tVApvzzJTRlLW40MEXb6K8vP
hEzJVD8+pRZmqzyEY4flezoVk/dS6LtL2OBFltfn1+daRgs6hmJyDiTrk/ZWx8DLs/iaPLUcZiC8
sbXkqHFAnJ5w8O9vhgYUal+2gTotrBl8FtGXePoAmV4hduPXgfNbbfyx/MDZexfkbs3i93osTviV
tDFxBoKZU6N9m4bOTpe6HMhIWsZEE7V4t81mYFI+i8Ue95xHyj80eBuuUG0QjqleYcpTF7c4bPUy
Eud01QF9awRJeyxuHXa5u/j48JyXYjJrQjl/Oqw76zI2+Cdfh3Ow3Z2HA7HMEkp8i3vSi4k7dpEK
lapXOcueIcYUh3QwaBfEUP2pAMvfyEXsEhF5JlxPuJ7JOF2oHH9Np47GgSxyzCmGuADOo7v1b4aM
VMoZApTVfeUD/aVcq0rk6o1NuDiG02Dn0iHwqLvn6K7vxXOnX4E7adNKzf/edrE3fXv/p66hnXdJ
LP3QTe6PVtfQjReM6HiBMYSq4pABBtCNcCNqYLW4bXoHO3bM1pHV7A27QFatpPfiTWHlbKpJIGdh
DK1JhIktXqdhOhQlXBudl55Jm1fatS4fjIkkLrl0O7ZmMDtOSmYCpiIVByibJcXSDLg+vPqHOzIO
N8znqPB5mej2PQPWPhVhvSWD4Q7FTAg6nb5+PGllk0joQUjihc05Wphz7Wr/G2SyD1y4pGk4v+3O
UJ55K/R+pKTDnJnVQHRlwgrnF7rzsghphPOxsLkbdQkKH4Q6EGbO8KExgA2tRQ92jfZVFCtyhqhf
r9PYzFFVXOvvmE6w6kUh/TM5l0fTrMaGjgUczKZ1P/XpMiSudso7jZYpPN2qwXUKJfTV0y0YmJQo
qN6rtm5HZyUjc6dA6pz8uD/WPWoTVTHX1mY16UMzHsw3HcUvIaxIuCPx+aFywQnE/40LCutRoEad
p/SC8WFAhSsiRjjl8jFIcH51P3MVczGFV4fqMwfzbq2h2aKxE1VbUJKzgS3/f8LiPMZEdNrOjGhs
QqWGtePc2FrYf8uIruMiLOZ7DYWxsjjbij20sVRyynxUklo0iD0eB9ZsorI9ShUTSnNx7AydnasE
PGONmUsb/06jIHyMSThB4opEr6otjp72EiILBqITMk4b9EuBm4Gm9S7IRRO/AS5KpKaofl8Wwwgd
aYJ5U/S/7LA4yYcT+uTVFtWL0iFjS2b3hIyuAX+G9dJOVCS9jU8/eFyQpt/wQ31vG5kbiP3VmEZ/
77HCD8tX8zGQhEg4oxZOU0QSviOZ9QDlQk23hcpb0vcrt5jO18vehj4w7f2su2qxt3K5wXsd/gIr
6nys2xPxo75Me7SLoot/V7MYJ941KM6hzoQszUFHzTZWpulMQnJERHp05MfqLj+faKcM6PhMfbjv
W922l7Kct6mgcjK7FYV5USzRugmxiHZYvAtWgMf7cVV2XkktLQa7seT57DVNfkLhEJd+MuJdmDR+
382CwbKDgVNjacuj5ZtUHdwdfCGPGYmDN2pTXHjY0kz/su7Ybw1I+nd9H7JRmSTQRyMsNk6OW7U3
EVmDPDX8j7fTlwRAjRHtmgzRswZuXKYPIaJO9n0JkcfWxCd6CPysBltLjH7qOMPSlBc1FqzNqLBk
lx0DSs11gD3RJwbTejcR5S/MnO5PSVi6k9URh2WCnd8LchKhQB/mKmbdA85lagqOZw6UOTgqpWBi
GD1oWS0iIpreZKiacUGU7yjtRiKHb4sdAV4LzerqJyQ2pAxqbvwlW6gbMMrcMa8mnKVexWIwO9bI
sNxtDJEgZHFM6kDuSzrbm3N75oV53CcQwuZRAAORQCu8hTg63YfLI6MRdmnzBrbnxB2zlcS1nMm5
YNGUIc0VOdwZ2OcXZy3ZsZqg3iZquZL4GSo/Zf88J0KkOn6TviWushi+WnDsDCJyLpgZorHvObhF
Rv7W5KNUbh0geuq5AmsSLsJkZqAWChQ3V65K3ZlRvMzAQEvoRCVxiHHoonGeb/RQw5wI4/SeFpDt
XEIh8eFqYm8DhnXhWmIR83yQ+Bg13oFe5oZSROsHZLD/poL6Od/0FeebUDUszogiCfonHiZ8CzDQ
3k7nA+dx3Y457HjRrm3SSu7dsY4InxLe1sDWdjzH0JKfMWKizb6FqJdaXAuq0ice+ezNN3H2m9Eq
yNxorE+hmMumXjhKJh5cyy1RpCaJ5V6xm//4WF3WFh5bYLrs//+YRTqtIjOOTvQhqDjZB3P7tlkV
rGcQnpJn+YjMQp9oLLPZIgaCkfhL0Gj4S8KOr2GenD3KE4Au6hGgYHIgY0mPe6/358fsTZ8RJtWi
H6sDH/jQStUNSpJVeE2fRv2yjRZIw6r9T8IQI0h8oW1qO4o9xaqB/T3yRFaW0rDjITqAdmhCzYNw
OCZOvUSqvZx3Y0W1C34kyvXdZLS8Ay8MBnaAjQ169zXU9hji8K/ENWzKkY9JWdAn3Hx88m9wVPYh
avCxybqkv2jgVgLfeq92tYcOyj1GVH0Kq9Rmg/IOpVZzjiYD5e5GAllOG3SROQAaRFC5ILWIE3dq
f1JxxQb1UkocpBISRk3WER9BoimXYZP9PecOoppjVM6rGSQs9XFN3F/t5IuRKBQs9IlFZTNsXei+
R+wDYy9YuxwE16kp8TTlqSohzxObFNmcH/BBXTE/exm5Wx/C0yhd0+saKD8H31mpoptPxj22AHXt
F1aY6O81UL8/96EssofETL2vOcdwnCQE1HYzRVnkb6RZVobz7E7n1nWqXs3aJ9osDKZhiZMD2sar
DZ8SR4sbulJbS3dgXUBhIzQCuKzkNr62FAtPMsHTKIR60w6ipTiBD3DzVGC9utFNZugmzrV4sCPc
n0/sUvwR1ulutF532gABQXZBITfueHCk1j08jaN4pem0LDAq5IbcHgeNL+Hy8q2xAoe48J1fBNiX
PYcjCV7+jwzehwcWoA7mZ8nXX1OC3JbajNoedYZu6+1pZ1lnwEJEoAHAAoCmq6F7RcVRU5PyD7m9
0hmnsXYvAICWlRBLXFnfRH8OzSMpxC+8WRvdOnNxQa+tv6PuHndhYeFQMXFXs4p6abp4vGXu6DxG
bx3ioUrt1e5unF4dx9rSgLQxh5HzK6PmbQee8wu0S1eZ2SEanh3qGwhpIxAT1oWTgjvA12FMRPDr
I3btnUv+w6Zq6KGnv4sswSl20/sWi6/fLCwxgHqNAfuR8FcwdNMYvBMPZ4SpyakPrxW1RKCLQvo4
x1luGxOkLYSclSQay6WUHlAjg84+XtQcI0FCOB1gGZ1/m2P6UQbkYrZeoVtPwwHzlYz6h98OLJCV
BDyhtCeS9wIKXnicLHCLJC3C4qkS6swChXDvf3WPWZh8hHcOHj+9iAdQbJbIaYV7qHnzARWZhOJZ
BfKJU8XxeTYaBgU+bv1t96AE1BfaOYbw9T1cdi+KsoA/f/9U3YeckQvp3OBoUXK1k/saRUkpyRIQ
PLelQi0rQHGwIOsEpMHbED6D8sWRJvf0Dm5L2IrxsDOqhtoWk2o4VkPZayPlh7wKWUskJlsO4Zv/
1X94ALdoqLccLzZRDUAVW2oDUsg/FtT70uj4gk2pJcjjiTbPpGaMH0kebUTjMRwweRIK6O13UQih
ZVtVeMh26AsPHLS5gf/GVvDgJLtv1VlZqhqvtUJ3YRGoJTVWIatWjSofCFAk8X03AMi81Feu7jBU
KT4Jmv8AGfs1ZKMLDDKOCxEGvDDrcKmo3YNvhl2xMK3otTpWeai3zrg0rcWmoqqUfgg887NbipYV
9evVQiwZc9VT8F6uhTASnBthlW5DJT7my+BfR19aqVgESzIn9tMhFJhTj3JVKTfEXR+Un3HfQAbI
6+mEsa9Rn2PF8F9lHJII3WzQbKw9Xp2Eo8dxRm31L8mXHsSlvMaVZGAhye0PRiUMHY3VYF/kGZXW
kDZH0D7Uim+mfFhM7T9M/qloIXevdW/f9sc6CwJ2SPXXhP6aC3mx9R/Pofcjnlet9Aa4coXBLjy0
SnTAY7cqPKnYST1CsCLmjwb3cej/istSlWG3v6TW2ikUCZiCV18W2mAjUyl+hYlsF4sTWOVRWfWa
7thFFBwm02Dzt2kFwJnNdLxZXKfEIjqR26ZFZFC6lKvxBAwUAdufTYHuHnBm/5C7mO4XdaDY36Nt
u+4jhnofZCNL68XtUEjI208Mcag+9fO+yS0pKS5IM0j5HdtLKrdrP9XlHOQigPm3nQwHQI9yK5dG
EFB3FooThsLOhVk9MexxjtwQV22SNUKTPYHNX0lKM/KUKiX/MneMrrN2CM1s2L/NjNRvLtyalrov
NvPBei18fICHXqMxZjJ3wD2f09mSTcOiebaEXFtlEOwapd9AGFuK5bebLuP0Eiase0YHnLL+RUDa
QOdL6KZ2gmExeyr2fxgcmBrGaihhURdnROaP/RRoPLwvyL6dVpbt/fAWqIC+hSwoXQjaCsi57+aN
PPh9hy25ogM8WzkHtdLmxNnQwTLflgYH5OJZ7KdUydYS6E04ZcCq46pYwRfcCeas9EsvxqECJt15
OTnVy3bGNwb0T95Ea60zEem/g92mTT1IbD+ZF57UgdFAKjbuAq6nr8SvxjyawH+8G4QzhL59+w/M
UaYClX2Rn7vsJNoZYIfkVGV+ZVH27ppRAYl7xPXzYL71nIXZf1pVKxWjo8113/RgBLmFw7kEjkoX
qxQYcDw/YbtN024h+vmgNobZtppmyrj/u9XD52hL5w2UiPDfALKrqV3GLidobTIOJ87+NNNrfZBY
pKwVwqTuzv5ZJasVked096p9FidRdu5KWt1/XjFPss3el2g0yndvU+Np6FjwUNYy3UdgSdtxhbP2
26j7/3nE97voFhO9Q4VIBa1zeHmFNADkFPnyj8thau68ECEK+8700iRrFsd8lU0ItAzDe21ON7tk
0ryZbwS/n9q0uLLb8oL8YcWlzh8WQzM2WDIez6afNUivN6b8GlviX7jIFS3MRylvFh9kdPW5x+8O
re0pwOeCmtKuIs6XkPy6HOWmRfcHNsMLK3i29GQZ1QV6gEjca64od3+OtDkiUr8bdMsPKPZVmC08
orteC2yRYjAOsR256l23DcpMQ2VHDNOOmcpNiP6ESCd3dTOuBmL1bQ+pdkF6Waxw0zoOnTKVZzSI
aIyasPZULobjq/JTgytCXiSmq+2oMjzSU+CpOuZVTH6und7Z6bQ3fikwj36CIBwynzoztMVu2l8s
tg3KTDun1aSBMvfd3jjzjW46CyaV8WBeaw8w9e3tMXIk24zSeFP8OieJsyJfsc9PvDJQQPAmkFUn
9y3dnwXQujNUI5WRvpmQfk+GAPCBjToJKcM6bsyQSTjYKZerktmAmVFVtRTSx0FTddQX3njWnDji
wfhcfwwMvRhQiW6w7bCXEPOxo7sxU9OD/677HpjpwTvsq6KZ4jpgNCAugx2eCuREHmqbchkvtYVO
TLFACFsAXzj/AQ5cZj8Qu0U8qyysx8NPSQvyqjtAqt7UhYq6pO99ksml5EuIMbCocQM1Ss9UqTQ9
NSTduCVaZSIIkhzOeTj2QKSjiMiSFJwfEYdGnvH2f1qUqsXpomIXVQjTc17GMbBeMuk+nrFHto+G
4LhYeI9PjgXvSXAtQevnUAapY4UVP1/Q1NDlROgeYei2G/8BZ0Hg6Bc6VlkUK9iziDg9YaSjFCMm
VCaH4pnzMOfjwJuTFhCfsfCXOxib6CGSkqZDF/jchHTaQpn9cS9wrOAzOPp79pmh3ectUwLJcRd4
T8Xn5OPV4wDl1rbWW4o+NSsMlvoVQLoCBr3d8hmLyMA/d2F7Jft8MUvjlBEr53xwYnrm+OlO+mWF
8kg0q+UhSqMfvbskioiE7M0bnt3IWUW7cw8Wrzpjh3Bhnf82Kc1E2vsRd0Ax7KXQfWoQlbrQnWmy
h7RKG3xAZzshPkrdfmKGMTYpNy3xCuUi2udx+1W4zCTXA3c8xnZd9Yt797aIONZCRtxb+UOddg+j
jxR4GBiNvWa2l6tIk2lD5gWWPNXzfF7UVKN/szbRFBQ+QPi6Fx68QvjrbArB01HWVPP/UHyipkEs
eYSxrfP4zVXNbyi+3kuCY1zcB6t++alxYG1eqUp8XQotog+uvftROpcV6lwICM3U2yqd5ncCTQiu
rW0nmdKu7i9/AVW5DQunC5DVB9xTKltvRhLWI0Pi1SBpsWNPxiR0b0mDSo4MzVV/AEVhPbsfP2bI
ZHzhcL9V0hsp9YHTDcv908dEMVgNz4zc5Emx9Dadb94slFNXgAtp77OWZm+X6Vv5sCE06GOR6Q+M
P1w5SgJh34AO8uVsjOD/gUNINluZIPYMjItto5ueU7WJ7Sdi88Cms6QrmolF/TwnNR+vSOGcP9Fr
Oo14tN3f+TFdSFfk1stHuIxw77ug/t10FwS4NAmgZgdN9fKEruIoad1X6fnkIRQdKLRbeUgfkE5o
Fns7UdYaO1mQ36y0MJ3+ftPz/ZTektOLVjU8GGONIWT76iO12afH0uTeQbTyH0BLKSAlw3j/gpDw
bS7oYmlEXQ6GKinPdOK/0OO1mtQqkyFJEncBQb8z9U1+CrrAg8odKyKM5TylE6TJUxcW7MEt641z
D53pcKglG1NejLpxhr31aPOtCGVr9GhtHBcOidNsiLGvJBHFfqiif5FiuhL6VV+pUwWBotloAvfI
/eiM0n4H6+Xj0Gk8pgOdD8J5JW2UNpgNZ4KqwSNV7IcI0VSDjYIpDlgOmE5hvVE4t5zfLyZrTHkB
MdKKmUyA3GUkkkuf5KmAPi6wSpx98DIxxqfg39Eh2Wm6cfIMj9qTdSQl4f0Cd7FTZv7Ec5vMkhyL
rC/jQ/uQ+mWTPrTCP771tXOfhZWsdIhtz60sEu8XWLVA7NVFbPkAMD9z4M17X1KfbTZlRYHDzUOk
hcqmeBvtiGJundn7Mp6lv50XAOqsoz9fu4gLQO8R/WcngT6Tj8YXRn46ZcYv0EAt2R67Do+se+U0
9seLRNUdZwTn2wrheVIlqSl7EcraVD9HIuWHzDL3RiFsB0nFGBZ9ggcgWhKjoxzLXfZ10kcP1NXM
yxvDd5CLTr0cJCK0GJqPoHUbP6jHXH6fGSIhNzbgsjikkcn8aDGgvLt0wuXzSvOkhZBhlknZwyEx
XeEmk4Sb4jAk+RqAl4vjpb+Cwd/ww1nRcYdK0PaWNDD5I3amip8pD2dkcOkUyImGk1wr8B93eB/v
IbE14cpo/fGclMWVEZSzgr3bmv6oEo2l3j9meQMOYpiQP0eFARH+OQlV5E1rIwNqaX5cIYkRqfD+
N8l77nBmEWS3L+aNpJP0odgH3GRE4fzf5d8AxebpF8BZcQ5sOqMifoeD8F8YMJ9y5JuDAwDfkT/N
GNewZHzM+Xwj0HggIMVH6e2LNlYtEY/QieexNlUruzcheBmxkqaCr0kiuDqPq0+wXMSzo0whQwEG
MCSAj8KfTohACvf8fbelHXHC+w+SMhKUh33QA2QdzTQzAVGB24GOrwjPYfN63aisOVil6zbNOm9K
+eCvOUxqZ9G2j2STlXeu+0oy2RUydnXkeoUh8C/N8GAN5/j/28yO6mWvqi9g9LwJKSwCWigiD6Mp
M/UruD3YQQ6PFhlkuYE2Z0g9gIFwHCqZwqMqG2pXp4TDeemUfjJskcj6BaiN5GuCyPmUCXUkIHmc
cOAbEch8ttnCItRfP3ERMDMffb4vOluUwPGPsG4UuoY+LHbory/AElXoGZAdIStBCTSZRegp9NiZ
enp5C3t4vLDiIvlIeX88pyZyzGe92XwOdZ16CZc8uZ2ojG1/kJRU9G5RN1AkJdZgNlvJAgnDK6/W
g7xKuA8rp+mPjEFHkg0q2DMD5M4W2Gd4UbJNsukOl7VU40/nM5UI1slmn4/dpvr+mxDrM20Nf+Tr
gDG6mJLGkJ7ubGhfaQ2R6+KtP7cA2Ni5S0w8TuJebW8gdUCUKNTSVJmlKmnJhjh/RQ5Uxy0VcZz+
3B8Odg/7ywDG3/5d9W+vFcFvJ3b1co6Hli1s7OFIfA4SilYZqEBvr06KdysjyJnBQWjRrR4zqgaM
P2Bw9TJf8XrHl27bp5GMxK8r29WKp04Doc2yzlybALJImvi9BIrObKwNtq0MAO27bij2VhIFsFkH
mYr2HqvFXsAsWss08G0MZ8vlFwTIAKtSXEjDdYbykzAzv4urxhjZ45z8rtPPyoXoVBNuLw33iHQX
e89kB10ZgSy3l6mdE+W5/nE9+6Z07agP7INQfEJ30WocZrL1YkiRUBlZPAX9ObgxJHFoUPLlygad
cDChREoEsw3Hs2JN908Wl35ToT4EfXSc34P1HN/E8D55VqnZoWlp1WMT/mxO1zaswwXL76T9qjhO
+LIrU2anEMywD41Pg5iyArloZOld7lhw5vihIS4Cu7RW+8IRsKATpQx5E5N14ojeZ8oQzfd0ONNk
FNHkDGlW6DYtDmb5Wf5ovcn1PVNwCkx/WxIyhfU2fkTupvHjch2wy/BEoLPw0UUj/lAU9sZ4DYAR
G4Vfo1e5P9LNMolClRWuTgqytk+q80t/xdm5lIEk7YpScwIwxOeqZHXQjz237fOwBUXxsZH3nfPz
VSDdW/kji+HqHTJBCfjctXYbxj4ab1qlVr6UGYkVp/+FqvpY5032Kc7tPD7rbTrjgseKK0G34mxY
2HqikZB2nqo9LUl3VD92OOoX4McKun978mUWSPA8u7Ye0SPYhiKFPfCuknGIP8t7r1KJJuh5Fxsq
ecLzfFWwpF2vif7u7QwXRD+rz8fozHUCmohTqBgBMJmA7fvUKdalg96eyUVdFwQL5Pyj8MlrZYG1
KtJZlHaOwugvZH1iYMzqN9YbzGoDhR6tByElOyX98gSfxRaIdJXoRSr70gEjiArDasf/blHEEby5
QX2ZZEWPUiZ/oBXZbQOa6nRj3glxGXqjJo7eFgtadCQmtaL0sYoj3v38XTYnk992ZJfwCkQY745V
o4RLwOygFGoH5pdLbqNFnEA1jbEMexs9ki5mcVjtLapYbqH9oIKlDJti8EAP2ocCVEeI6YOlSFsn
ClJqIsq0kZRE+KLd4+u0j3AYXv2aIgSuvmr0ZipJxAFrqvnqEMn+/YQgIHT1Q8EIozgSSrjGqhAl
t5YZ00Xbj+OEtpSsraTa0K4AT6tADdtnsKq+Gguswq9A4swJJKbWBxWdQWgDKnezCrIXnC84ulFP
05jYnQ7ZpMMaqBzA14658LZV4BG7P9NgfH+F/o2rZV4ZA4uiENInWqimVfM/bqNl2kdlKyj8PkcP
2Tiqt36Q0Y6mbVvyq2PUw3ZWJ8d44UPymcpFQ0ScyIv/ucUp7gzCgw5LwSo5//yDTeBd++KS7lE5
Re90Dk0PBm2/T92Aqw0zKxzci8NQVtrLgrmQZ44m2ng8fBx8f8vCZ/NC8SwVYp2tZ1BL8aBGmxJ6
xB8gJU7fh99bUZQp5JdqwrRqZApy4lqJqUwNk6qC9VmvWe/5d55PDBrdvferMniNo+/8epRJZqGe
0gUxt7SPrcrQcy/rDpMmLVy2QBOByWt2Yw8WSEt+MCrzE9zw7LeZDGdShfUzq4A3Ma+29K5J0/Z0
gF1k+YcWCLXlNmq51xnVqLNeNhbgrAh/h1nF7WFC19kHJcdNbP+DZWTe8y8gEOcpW0c0sMyiH3cF
EnjLZzLyyvtvN1g1qRWungZWf5OL0foO2JuKW4bsCGj8zYb7g4Knavrh4MEHGZ8twuXAVnX2kD82
s2trhyQv3ATPRaL13jZ59ssVK+qp0txQs1tugyDKkOfanlI+1DqyT9UZR4kMraiDxvh0FEO4DZQR
TAOKGuR/HTxNCSHzukOnUn0FWnLVi02U1bidrDzNf5Ilf51BpZopSflD1gWDwnguNX6zI7FUGkv2
CxUZRjgjSV2h8SG0wd3NXRLYWpIH34vA6Xjm7xVm3jIzwGFDkNHC4+VqakoNbMVUP5c3k9wCZmRE
TcxJMysZD4djwxPmsJo1IOtun6U2pPo6KrpkgiCyf2Ji01liEU01a/ZBuASKTUqIhF4gzk3G/f6Z
NwXD8OEOBT6lEYaDD3NisRXIVIbJsR7ybE9h41FXcFPzxE6EWlsrgtmW1ZjAu9Ark0y5ZsLZRADK
lwu9O0hAC99wvMnmp4c/NkxbGs4p5smjXlYDBWTLHfDjtAXrhGD0VXi5OAdxCUHkiNiqDai4pzj5
fmGJvOVAd23ZvnwAe5iwVwveE2Vfj7rjXS/zV9DRS+xFVz7ITSPfA13Jp1DQegr9a4e/7OA1tequ
9hGTOIT5w5LGbh5Qv3GZ5zWbmzZNPM5GIJpnUhlvImh5LtX+cleSZNbrLxdTbYV1+CiPYeWr/1Ca
Z3z/iH0EW0OhNN0FH5O3X9sd51u9rYXsbGrTG630gEygHN3ZPy/ypsQ/j4A8duA8JuKUhv23EDl/
yWh+t+E876NL3tT9zJPTHMQ3C910UHdDFhO5InGBFDzpbqbXBbAVFooqS9Qj+L4WaU8KySlas7wF
XoSdviBe2FqPCJvR4wfBICeUyv3Qe86vqb2DR7bQ7HoSk+uIS/Bg9+ybgoyj4nTW7myfvXZvNT6v
xOgTYcjk3pkxxmg6NYtAkumm2m0HTm6UywxXfV5twJYjzksan+SrRSbCKnMdFQtbeUuhOKSqIEqG
aogRbRA/QTKbngIcoHtenwqG7clJl0PHxkZaTbpV0vkIX/FMiSevQMyJI38y2wU2GElAfJmZ4sSX
hVFVqY4VFBN05Xkpu2rbjcRISRxYnbugssRnG3iuShawQVxfk0RcjUIuUNBEANa7Sg6DN0RNGugE
5bDUAElQ1YacGu/0c9qpp/ps4Tj7qlWHRvBHMkHyD6lDThSAN+cIXtiMaKUGBEEHWdi3JsQf+mEO
xUCCMsQv98lS6Y+AI0H0EY35HBfBzR3/CQLqlFN35zObMX0D1NTI8IKhaLUZwEgiXarj09vW1YVQ
fZffwY8E8JIdYSdlvLFIffQT/53Y5uSYjOWAecMlkleJTBKQLPjG4tqOwYzJmnL/tGUJ8xVJMQRA
cXFOL5HkdwNGfUIPzORoCpSP+MuL23ecm/DGvMFnACjGYoDEaEA/cKQJhrCNot49j4GbWl4XlZTF
wukFGhLyjyQc2NBMLlH2aruBS0IY8wRY6O8IjqilkJi2pz8DGzPpKJaA0JyOTtzRX5ABS3gxRJOn
7N/mgk0R2NODcVY1ith3/vmXb51OLv6XK0NGMFpVBIk+cC5jQ/dchv2T7a8zmnVEptZuPl3/TSH/
7Y3lHjX6M3a3AJOQ4sRlNJYs/IJ4L9Xi9ftb2a/J8zBU5OjgFoEf7LFSM/8AjxLsLsIFMN5p0d/0
pEFuCP2fojaC//YPA77Kywfo004/voVpEa5YFxDOQR/IJGNCkk6bi8ZZx9495RUTZJRHhSeFr6uY
uTB76X6TM9C6yZMV6dzZ3vOh5KHuaPNbeQ9PlxbGHO4ubcl+tuWzm9P3w5edBJheQbttZJoHOlZj
IPlcNNKPXuzWwETHFrgeB16IvmlqCHODZN1Ie5cnxKBMf4sWWmIOX1ijJZneVYywZunsVj32akiM
HhfRebMbwf/c+SdLQPigLerFWumRFXJZsFtssHu/YT0GAF8cXzJiY2X+B1s742jWYpHLaKfueeaw
GI8nAeQMH48XyNwKLJ2bw+ZwCtUTvBWFE5ziM1unXMBl2toFA3Dc5C5Xby2jraI/aT/ToDmdc3OL
qhuJgDvCRYlRCavOT/kNdCj4L+e5aK+TPp4uoCVzQNuN9W0sQoZ0sanRE6S+gJE8O/j0QLYREV5x
AO7jIYLnbMVi31W/oi5Nl2hxEw5Ao+1luG7BoeKpr7Agb1a26iXbXx98UpieYUvKIejYDc2s+wjv
SxPBzV+mX9Zr0fI5VLZVu+cMU8ugCxboxivmq0HxtcpYn1kA+ro8LOnBJKXxpcEEmWjgZJSe8nmO
KAp9oIOWLwtZ+q9r7OiAjbEuWtlsqkdpzOg3UC5wcdsH5sHoIjqj1RNJQeaxLKMAr8s9mDZCFIP0
xSLsEu0+7U1Z1y1FrDXt3n0+HgTDwjzGSLsSYu/cEzp9KAdKxUIeYIsKRy4S9vU5XGEeI9e4lWp+
xzTjkueF5f8+70ClI1kjB6RvOvd7H+E2fqw0FCi0Ud1cggiPVRtT28FP52YWltNAbg82JjP4alLK
9Apf9t9UMEIsNywZ5HZ1X4RQwRjADgSpRdEp3njGw9tk6OlkHzjC5VJJy1Vut2aMMTqf0yFaHqoz
PCoP2c9XJYQQnZcwXK+i/g0mwVm7yGusISOnpGiupqd484Jky4mQGzNOzItgv3SMYsI4YjHItV82
DhnP6hzp78uyHG7ECFRkPN5Vay8PPnjrFSeHBSSJTXk4UeEBnY50RFrLrammD5ZojA2LlmxpMnYp
5hMV96tBqwAzOg6irfH/6VvGCRu2bWSH3hd6BL6/8nfHU872Y6XGqKp6FtJ5cZUjLDFQpvg071el
zQqglFKLWJ8UjsSqhNQDNla8eXuKt+stWYROp8uYTnmOfMR2qzqXqMIfC593Ap0+fcXbTDGO0d84
Mfr23l65errTGI2WFoPegGWR9CMA5wGJxD8Wt264iEQcdVo951frEPCxRJkbJVyZHxww2yDVgj/r
sLLmZDWT8AOs2QHkyz/WdPfP0rcsG/HmnMRzfDpBsojp/uf9k4lz+IynJZn5qGYJZJVV76iO7Oli
izwUtdxBLTdlAvmV43ZtNqUJdcDWW7wiS4QT1OyyN0BfV1H56FtSMqMh3z0t0QFMBX3MUnqE8AyQ
2/q88SQwOPF3zGq2e8VgPJQoVOJ/UeLR+3qX6hg4vDkairEFWHylSfNfIgwtruJYB/9CapL0Q/BD
+R8YmkSEXJzHkrxh3fkrtsNhGMwQORavAh9Y7hjJfIgjw0QHeAuKiE7NuyB8us+YRbTE7vZK4fCX
zkwjZSHhk8Tue3ryCMXIMUb5kbF4KImk0LkP7c6xDVOrezG4uf+C2TjMWf3eEWteucG+8TWVrUQ1
BCYS4O1fc3zzIjXw5FmkKsNFen4Fbio089ChZuqLCoTOiEB53T1MWuL6SU2Uk6BPnti1mIRnV6xv
GAMMcjjYfhMXmcbmodbtj5kDoFzEODhIgXaNkdOi8SAkwOBRQno3ZS8VpqknPnJZcClWcj4eyaEB
Wjqtec59+ClD3oMdHFRvMxcVOgIi4gG295/JD95Mf+2nteEAQwOMuSM+i1D/Igd3cLiWCQJK3JYj
WI+D0TvuuuZEqhD95sygptXPmWziiMXlWtpfx3hmO7EEu1NLN1HMON0aoQhEAbMBdEcpSptn1v+j
SOJo8Q9BHZEEnWvyDNb0X+c1SHaZ5z8qeRfJutLFf0FM8i21826Nq2aEey9XKKioRao+m5tHPlbu
CtV+sn8GOknpnEX0CLdqL+WcLwWO38j+ndCKfQEb61+EO7FIKNMK9Ba2Re7Scj2IM0qUCRZ2JN4/
b1EBy0jlbFl5KXNWiXo0k6wzBHrZwaA4iWSiSOPUkV9kPODy+h6FgtyIVcGbClwum9k6+FZEHKWS
HTZPjXnROWMc+PwkUTM8KRZphCI2Yu+LB0nIoeKRuSeDNqaFOU55/guBmZYXfF/QlUCHvyz6dSAM
use4QP2R/nMooBtNpetJTfx9+kXy+k0lksdnM4V7yFNE7JBDexbDwNDrHnhsZs4YcE8qUjhn3/kU
pfnzatl55Jl2ciMPAJQEMSVOALBpfK+vSZhvR/sunkVVDmHNrTGgD2h636E7oiaPBgFDs1W5eQsb
lC/oJ3SgA5YmH2c3XY2XkqhTO5ZphHxbEpuAc6OIKrKe13mvdQDRabvidaekTjrbGDwA7c4jjx2V
z7/0wcUbOmtGYoP0EC2/iquept1mjf/X4chLiuAhWPFeecoAQzZiHhB3uyAA0EE+59fjO0S9FsTz
MlhlvZ7UrJgjYCKSz0m9ncSFmdQdmAr4CW8kQ3bePwzMJ4c15ZaMj2DACXodexTkKgcM5sUG9/Yi
zbWD47qFWL77HOCBbA8K2yAn2+5VbR/G3jCAkQH6Qom0GDosXqtwEQlXnAsYNs0Js2+yKgybD61C
88JxM6qa0yhmLWB9jmsOcz+1ma+g/Y8eVVZzyngt2C+000Aam+Wc2mRFJdi5JBB3ywuShmJ9amrT
EXo6nusKRiPdH/5j/Qh2BMscDCJss7XYbm85XooQlVgOhv41Fu56JwF4MdlWXMbiBdimu1VHON4U
/+un2N5iG84FomUQqM51g8g64FMusj0vHiGntavQADLBhPlX6yooaCrjn3DzHrkhv+QAVEsb6V8D
tKI8PGR4AVjuTMsSrJtd6Sfx3VTSE5FwZFFALhm9Zkzcm1PuebKOMW27hfHG20JtpuImzsyVRoXJ
nSeCfAnCuCydmyRhrkXHhnUIyev2rkxAMCJ3KURjJWtknjG6C47Av7UvC+HQqWAdTCq1lAXFtL7J
puectRGHwS3c8nkmevpEWBprHKDMLAVDxcexbfkmKgEoQ2pSZx9lv1fc/Djaq5UKeADxzq52945a
olCnEnF9RU6/qaRXIuQIWUC3VY87ObXw1QAoquU6IM2DyQSdWDHEQ+Mw4QycMPW3MMytXaYUalsv
ywwmoFM3yeY5P7YJkmGt795VXziuZV6GEkO7I+OuZ7Xk02HOhbgwnDNPzhaNVTyCLGZkXeQkEBjq
qI0ke+ptkVpKH/C+5FTqaeiKg6u4Jtk1HQBvuTXhoOmkX7J8vJFbF5+RyPbduPSzEiIzeUtUDLDz
Su7tyYgIEcS25uw9VSPUL9DM3WHtABlIbzltHtJpqVZgFRqN5HjGH/+vadclmYea+LLmYLlkqzbQ
64cBgOi39DhFuXiek4zYZjtqdwagMgPKR7rffIbh6MTGAj71Ae+1DvxP0sL2r/teayepzJ18UlUR
WTB6HAdm5HNlkpg8ceMBbThNVQhk6Akrkxjc3HGlPRJQRo+nzhTT1cRITRiKRamE/X0E1Z3lkf1c
81kmqxva7mZ+uITh+nng5MRV/atnJHhFNbvh7Cw4GoSWx3OH8wD62OoYp5sfiYXpFwLRTHJE8xiy
bt1Xdj/boz3J/SQP7FYZcJl8X/AQ5s8XE/4fgeNx5BVygOFUyGvNO6++GXcWmxfb+eCdaYj8Q7/1
rrb+Dvqehxtf6fWtunzH6eOKX7mZGws0fcbXTJxUBTGolCVwWJ7+mVsmmGb/Atys/QQyboRb5X+7
Q16vgT9N433JB11hIDkTAyL8UOfcc2PjqfjzPbzVOuBnSR/jH3nrM9iTwjcv1qNrxP8Jw9oPi7yG
u4aT9vidaSVfPLxNzHD78o8UTVSTTWeTwMmau1CsLiENzbT+wifRT8HzdQ5K1/aCxKRIwBqCm2+c
8XrMXyXILBzh7bYKNmusKrX5DnCXAwbUvNuedz/YaPRp6MjO2vOMoJp7TcI50SsJyWeL1ab80VVq
zymk3xstIeuGZyG2OWgLXyq9DGm8QBv1yTleBz7eLip1k0Dd68Mx9m3dCMdjyyvXEwOpsEJfNrlv
ToIRpav7iAt0vbXtYoaYZtFxCuVLx7oR+zGHmrTImHmRCbz72p+WXI4Rzq4eY5Dfl/h2R1dvKSQ2
JYk0phDUzYuE+P5S0aEXQoctM81c+plck4UTkrI1+tWciLbOX0+99QhBaqduxfmoWfqY3diclHgw
ofw0lCtR91kGOuFPtSXj33Qs/XiQsP36U0yJUb14P44WwnX+Gz7ibuPz98JG/wKPihAakThX14sU
egacCe1qmjIywsjdgOg0F877tTqm4RIVVf3rfZHHZxTNUdwvpLYvbDNPWt8NXXKuAi+xBYt22XDD
3kGzlIe6PuGmay7pDSPXccM+dnkQKR15pAqkqrzKHxd5Wt8A8YyOiH7EDmYMDlgcXHP8MwLCgxtG
h05cdOs6MNlyocHrwgqdE/mKzqSV6ivQIOHnDnl8xTKIsj7Ivl14zWUYmS5M7ng6JuT/9zZncoh/
tkNArVtYdZAWCwWoUhv6AbFTaE3PptkoVDcRWku188HFVBSfzPjcrVNyQBiDJj4VxMIl+eI5d9z+
mgv1OFqpGti2TV2d3udpLA8q7hRVXjCjsR5gZ7RMXrmRW2Do+qmkosixaQRnwEpkVBBwsOz2Iihx
NLf79n6KvQ5C1s7/ldRLi+sAx/YujzlHBSijYZEZr2CgMEy8/pQXcSfG3TDai6Bypm2AEtKYOifH
r429eeKbiNs+N8Ilp6C1ruJXa1Q433JODCx70lLqlq/gy+PyEo1+lFSSfRtX/su8uW+8FelI/wfc
LdTEXcddG4ZVv7S5jUBSFBEKYnz90zO+EmuHi6mdaeATC4pTG5A+GQwbpKgvbm+TYXlDR8cCHiTh
XNYaclF/Arsv4Z7Om49poXXmOF4Iy7n0mq/q/QeaehahX7fPhiDD1YqqVc+roq3m8DXCPIutaYHC
Qku/61yY2qVvJ5wKuPGafDBz+UuEmmWHfHKCgYsUSayOrPFZPq1LHx64dlvFXU6rEgdn/E2OLip6
dCbe0nV4qH6LtPXzXz239H6IKjDUZIJK3tUJVW++TMIRT9/DdStOV8DqO3ACIyNUO5QKwN4Qlkv8
y18gaspGM3dfc0xUxhikpvhyyCHJBmoD/s2yBEEbYyTuLEtzf40sKgbFC5K/gC7Wj+N9iak6jx3G
ZKlp40NtZq17JwW/BsnWvQXbO6VbFIVx54uxqwGn2p56mCKvkZQCkcIE6W6DCiJH7PQcjiQtzADe
isWcy2Y+evStGmkADob4SwOtgMh5O4iOrMFWlWJsHW8yOgzqKGKms9m7RUKKWoPKPclPe4+kEHfN
HKw8hOtN1HaoHdTsSMJN0vu5w4Ut5QeP4goGS8uT1aTHz3FgNVscU3kMa9fLWdCSjUsUBP0FF7yR
Np0cSUPvHOJNIeDplnKwDPfxb09o5neDd1kRhuZUpUg7ynJedKB5ryW8VVbxURuHB20ziO2z5rzj
Z2WrfkSAxQzrbGx3JsZjQpCW6ZT0OqmFlgJlrESquFi3D50+YzI6v1WPjBI90ja9Cb8Zx96XL8cC
f3y/BvQPv8Smddq/b/ZAfw0q4ycmuKd9F2bZ0KCdpeL2AGKvTISp3KoO0GFWhSHi5q3uOuPtKNtu
rWrpY2Yue6muN9EMAJC6QRu8d0720JDQbZgQvCR4M6sCODiNLsS8fq2oQ2pMyz4afGFcg3jAXivU
woXwMOijN5NVNAnE+ZT8/QY/JML/m3pQ+YST9ijQ8uFkj6/s2HXpdSZo20Li+sh3Vmk9/fRM6IkU
36Wj1joPJNyCOq/425vWEzj3pZeMXTOf4WtyYdbvwQiZsLFl107FYlO2Fli+hfWICmX1mOsaARqs
gIapLq2Xr+AXri+VfeJ7X+3W97BUaNm+lLfqxoGR7aY5mj/hyLImAgDmhW3y+4pV3yfw+aAktKA2
MdSLjSAi5AZRzU2umn1vdGxfWjXuVPeEg//85nJOsXAATQOEcIBDlUfhElmBlVoPDuNoRcqkDpOS
DQg9UEHPbSZR9XFjd3FrIarj8uKIb+CX0RyKsAoo2tNNILuqpi2Sk8RobPmaOpOTS1LVevo64ubJ
NBt9eerIPk4OsFE/33/G4pfGyDU9QFFCa9jxy5YtIKo/2M2N73lg9k+iIv6X0YLdZMMSAw3EM6Pa
2P8KKgyk78DWr1q5eXj3qGf4gwByvIFsc9PadMmZt0xQmd1nzSVUT1i34W8NMTcHoUuR2bQKVfpy
nKU8RS7p0rWw7FEqQ5q1146+qayuFmlkb1hHScdXVzEIhOm/R6D0KcwjnYw0KOfmDlYOHLdadbuS
2Vdl5SsspBiOZAREQWz9rkyBRu2lHGNYGHgtxykhwhpkcpMWX40+NYn2jIDvg/6z94m8yfW6iiKq
FqzAKsXrvO3VMRdL9GAxa6qMgvqWZmo6b7NbIqyUZfWILUZmdyawzEz2ATgLiIAVfDHWklnwT63W
3pWzaNcSYmeJe9QIEVeqytPcW2ErSpfXHflJLJjfC6iXklnoWejKiu9BCkFx1ij1fmibOIDYUaiF
OZAI4B7CWdXYbnBU80xqXYkyvKEZbJQ5Zrc/UNY1C1o8jJGNoLTZMKbZ0F7ZCFIIF0NxaqnGeqRm
3zcxHLpT5iuUoiqm+leLZpe2IFYdgmlBcne0ots7loTTf0AaX4FOCYRn05d7RBbfzwQ5n5B+5xwu
EpF5sxQaEsuj9MWmb7zIihi3++DSLi8eKIHJzgQpATtNIVaEn90xeEZHzIBMYFrYc695j9wT5RPz
MoFBysPMPcVvKflRECsyetEkJ8nFIs9069RxjBssSUMDthB0v4OEVg7W3J2uqzXIhnCXc53IcSHB
JlGOXuBOo5BxXKm7exzYAAjJYj1IVU2RXPfTN8ejc+E9WmQzPBR9SJ5MiCIP2A7y9Cny/UiZsH0W
ZCgbQ9LchhrxTlIwV7q+ME531BF67rqImgagweaf5HeYqf4yez6lXAH6+08DBDaTERT06Urce/MR
/BYSfQJZ64u5Eg4DA2DFcF3hdMc02K7aDg084+P52KcwIChSMkOsPfRnuk7CuVDqE1n67x++sexr
FuwR15Gqnu7QwFDSHadbYpflOXbZCanXcJIIbrb4oEBRaA77x/LOe/G2CkrL/XPXq5iqMbrZFl3C
gQRsOyz+54GOUV0AY9t8x5IhF7Q5eYWFsvpaU+BlSB4e29HScIQrtpMREMet8JnUfgyFYsToqbPv
hM65flV0pkynlxYaEAoRv3YU2YPUZqHAPbRBsJ8PxbrVGE63PLbqN5G+Jl+GhqSBavReVLKRngBq
fEDGyctIWuREE60qjYQ+iP9s54DQ5zOYuuLhBk7OGSuEIHRTxSgf6OIMtvPyIEj78ePREjQOuJv/
3D6obcu7YTfXq1ZIQ1jJ/ZylBWpfUm9dogo6k78L0TDrMAizJzBev4FudBoBKFclvwoELsDco+Em
f3MZAzzFcE3LQfwr3B4IcambQ/ZDkfIfCk4X0mbl8R2BXuXMcQYCvHV8U8f6gbrmAc7XpaVguYOC
UjXnIothHlbltMXtaKUNelcfAl9NVU1DddEEN1oP95kgJxHjQasIQgwZaVeKY0akr2wYMlsvkjMM
klMT31rrOcrpOuX6ThBRBpP1HwFWHIkSm1293rVVaIVkiXQwdROjP4l4db8FLBxLQiCLYvKLoN+u
vo43+O1tFIKSmaAodTeeka5tLRqcTDu+qXeOHLgMNOsLmNOojNUwFa6NpKGN1giVdNsDzvjHyypV
6UBDo/l3cw9qRYo7PWPK9UlCR1McXIhsFiM2/HO2JaI5WKJtL+aCuK+G2niV0ImmoEvytyV6kYsQ
Fj7jnFBzFwAn5WGrX00eVVZ4q8XKeQoGUIerXAFHoaEiD1JshXXHOnlJJRmZVDocCOfcfjnM+L8D
TlnoRj7o3zJ0Lx1ZkaxU/GFkEc2NigdxrAQJeXapk44MeApRkEy37ai/Dw+81c73mU18LCymZe9C
iH2enoFF4SVzNaHF4BXwUZlFCUPQL9lcXpOJTl8/yMJkj2lXMypylETB4GsMITYRnmrvB3y7+Sko
Zxsk5fkiGuWqAtUbMjw9YEzbyCHjDj9VbQ6lhep3OkHmtIEw3m41JMDmFpSTAyU8ejfWoR50IrPK
F13IlkBBrR1yajZLZMrUitUmOVP4dqZpu0bhk4l2VyX7fsWadD/srt+e3yWkPir0R5EKhvgI1e1U
nbROtbnDOj3i4RnoTlI9Zl/A4Hp1wK+odCKiUw3qbECrSA2kEZhDBIqUQlvasmNsNfcj8IHguA3C
2illNjD4w6p+Kmifu6dMp5DHYnqDYO7D++iOQnfcRBpqEJMBRg8ntPc2M/FR8Wbp1oBI/uckA/La
R32MlGy4ygaYbGpnQPi4sOG8A67U10/pQeoyD6B2F9tPtg9ct69ASpcarLLZO6vNeZFnmmIfRTxV
UCAW7fzodcGR7qUrqT3Hw12vPyxfQcC3fLVHg1Jv7vMfsvhyLu14TzIsFU0425GuMvOJ7+hxw/9w
LyEno/w4nW+Nip9JMimEqmV9nV8l/4jt2FfAFGIM/54J2YviUPQ+Dmzh7isVzzlNco5HacCyBCR9
TWl6Ou+38tLquOT5j+5w7g+Wy47kl+WSwiKAzzK9r1/t9eaAQ4JYGbGvKqvkF079ChKXNjTM9Dxj
clKgYSE7sJMH7vuUdrdCLC9LXnIZvgCQ5gecORyimapT2JjYF/9cA3DPVH0BBOBaI7qXgAKY85He
0QSGGHcJY+iFhh5uhoHxiDS1t7tJ4MYaYwbJZu6e+cI6b8B06rD++6kyUUluSv7pkvcMIpEyQvr3
1Tkcme4mvI4tH79ka9CZOsL1nbJgJR8ral9HcWfibJfpo/DhaTj92FZqsNwJf+jkHEhOGVSTzM/k
7/oYA8THPqDufd3iNXXj+kU4IJ05hOvT+p0/eYL4q8wzqKNINHyGPmpkJ7Iyz/qKiDLvb9g6JTYH
IE4X0qnhkOs6OWHNWDqs24CWCggMkaQSsWrAc0W4SGrx9tIn5JoKMYYyrk09TNkvH02SRate1KXQ
ehss29KpSJGgg1mYHre2Rh2T9rqQs09ACe7Q+qs6gEERS0VV5k+DpTjscUOHTA0+5CLIR9b+asPQ
GZqw1anqxt02TRfpJCOQiRMOYYnsZketdVQyOv85fq/02Tr053vZKOTvWw==
`protect end_protected
